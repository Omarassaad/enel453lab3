library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	8113	)	,
(	8090	)	,
(	8068	)	,
(	8046	)	,
(	8024	)	,
(	8001	)	,
(	7979	)	,
(	7957	)	,
(	7935	)	,
(	7914	)	,
(	7892	)	,
(	7870	)	,
(	7848	)	,
(	7827	)	,
(	7805	)	,
(	7783	)	,
(	7762	)	,
(	7741	)	,
(	7719	)	,
(	7698	)	,
(	7677	)	,
(	7655	)	,
(	7634	)	,
(	7613	)	,
(	7592	)	,
(	7571	)	,
(	7550	)	,
(	7530	)	,
(	7509	)	,
(	7488	)	,
(	7467	)	,
(	7447	)	,
(	7426	)	,
(	7406	)	,
(	7385	)	,
(	7365	)	,
(	7345	)	,
(	7324	)	,
(	7304	)	,
(	7284	)	,
(	7264	)	,
(	7244	)	,
(	7224	)	,
(	7204	)	,
(	7184	)	,
(	7164	)	,
(	7144	)	,
(	7124	)	,
(	7105	)	,
(	7085	)	,
(	7066	)	,
(	7046	)	,
(	7027	)	,
(	7007	)	,
(	6988	)	,
(	6968	)	,
(	6949	)	,
(	6930	)	,
(	6911	)	,
(	6892	)	,
(	6873	)	,
(	6854	)	,
(	6835	)	,
(	6816	)	,
(	6797	)	,
(	6778	)	,
(	6760	)	,
(	6741	)	,
(	6722	)	,
(	6704	)	,
(	6685	)	,
(	6667	)	,
(	6648	)	,
(	6630	)	,
(	6612	)	,
(	6594	)	,
(	6575	)	,
(	6557	)	,
(	6539	)	,
(	6521	)	,
(	6503	)	,
(	6485	)	,
(	6467	)	,
(	6449	)	,
(	6432	)	,
(	6414	)	,
(	6396	)	,
(	6379	)	,
(	6361	)	,
(	6343	)	,
(	6326	)	,
(	6308	)	,
(	6291	)	,
(	6274	)	,
(	6256	)	,
(	6239	)	,
(	6222	)	,
(	6205	)	,
(	6188	)	,
(	6171	)	,
(	6154	)	,
(	6137	)	,
(	6120	)	,
(	6103	)	,
(	6086	)	,
(	6069	)	,
(	6053	)	,
(	6036	)	,
(	6019	)	,
(	6003	)	,
(	5986	)	,
(	5970	)	,
(	5954	)	,
(	5937	)	,
(	5921	)	,
(	5905	)	,
(	5888	)	,
(	5872	)	,
(	5856	)	,
(	5840	)	,
(	5824	)	,
(	5808	)	,
(	5792	)	,
(	5776	)	,
(	5760	)	,
(	5744	)	,
(	5729	)	,
(	5713	)	,
(	5697	)	,
(	5682	)	,
(	5666	)	,
(	5650	)	,
(	5635	)	,
(	5620	)	,
(	5604	)	,
(	5589	)	,
(	5574	)	,
(	5558	)	,
(	5543	)	,
(	5528	)	,
(	5513	)	,
(	5498	)	,
(	5483	)	,
(	5468	)	,
(	5453	)	,
(	5438	)	,
(	5423	)	,
(	5408	)	,
(	5393	)	,
(	5379	)	,
(	5364	)	,
(	5349	)	,
(	5335	)	,
(	5320	)	,
(	5306	)	,
(	5291	)	,
(	5277	)	,
(	5262	)	,
(	5248	)	,
(	5234	)	,
(	5220	)	,
(	5205	)	,
(	5191	)	,
(	5177	)	,
(	5163	)	,
(	5149	)	,
(	5135	)	,
(	5121	)	,
(	5107	)	,
(	5093	)	,
(	5079	)	,
(	5066	)	,
(	5052	)	,
(	5038	)	,
(	5025	)	,
(	5011	)	,
(	4997	)	,
(	4984	)	,
(	4970	)	,
(	4957	)	,
(	4943	)	,
(	4930	)	,
(	4917	)	,
(	4904	)	,
(	4890	)	,
(	4877	)	,
(	4864	)	,
(	4851	)	,
(	4838	)	,
(	4825	)	,
(	4812	)	,
(	4799	)	,
(	4786	)	,
(	4773	)	,
(	4760	)	,
(	4747	)	,
(	4734	)	,
(	4722	)	,
(	4709	)	,
(	4696	)	,
(	4684	)	,
(	4671	)	,
(	4659	)	,
(	4646	)	,
(	4634	)	,
(	4621	)	,
(	4609	)	,
(	4597	)	,
(	4584	)	,
(	4572	)	,
(	4560	)	,
(	4548	)	,
(	4536	)	,
(	4524	)	,
(	4511	)	,
(	4499	)	,
(	4487	)	,
(	4475	)	,
(	4464	)	,
(	4452	)	,
(	4440	)	,
(	4428	)	,
(	4416	)	,
(	4405	)	,
(	4393	)	,
(	4381	)	,
(	4370	)	,
(	4358	)	,
(	4346	)	,
(	4335	)	,
(	4323	)	,
(	4312	)	,
(	4301	)	,
(	4289	)	,
(	4278	)	,
(	4267	)	,
(	4255	)	,
(	4244	)	,
(	4233	)	,
(	4222	)	,
(	4211	)	,
(	4200	)	,
(	4189	)	,
(	4178	)	,
(	4167	)	,
(	4156	)	,
(	4145	)	,
(	4134	)	,
(	4123	)	,
(	4112	)	,
(	4102	)	,
(	4091	)	,
(	4080	)	,
(	4070	)	,
(	4059	)	,
(	4048	)	,
(	4038	)	,
(	4027	)	,
(	4017	)	,
(	4006	)	,
(	3996	)	,
(	3986	)	,
(	3975	)	,
(	3965	)	,
(	3955	)	,
(	3944	)	,
(	3934	)	,
(	3924	)	,
(	3914	)	,
(	3904	)	,
(	3894	)	,
(	3884	)	,
(	3874	)	,
(	3864	)	,
(	3854	)	,
(	3844	)	,
(	3834	)	,
(	3824	)	,
(	3814	)	,
(	3804	)	,
(	3795	)	,
(	3785	)	,
(	3775	)	,
(	3766	)	,
(	3756	)	,
(	3746	)	,
(	3737	)	,
(	3727	)	,
(	3718	)	,
(	3708	)	,
(	3699	)	,
(	3689	)	,
(	3680	)	,
(	3671	)	,
(	3661	)	,
(	3652	)	,
(	3643	)	,
(	3634	)	,
(	3624	)	,
(	3615	)	,
(	3606	)	,
(	3597	)	,
(	3588	)	,
(	3579	)	,
(	3570	)	,
(	3561	)	,
(	3552	)	,
(	3543	)	,
(	3534	)	,
(	3525	)	,
(	3517	)	,
(	3508	)	,
(	3499	)	,
(	3490	)	,
(	3482	)	,
(	3473	)	,
(	3464	)	,
(	3456	)	,
(	3447	)	,
(	3438	)	,
(	3430	)	,
(	3421	)	,
(	3413	)	,
(	3405	)	,
(	3396	)	,
(	3388	)	,
(	3379	)	,
(	3371	)	,
(	3363	)	,
(	3354	)	,
(	3346	)	,
(	3338	)	,
(	3330	)	,
(	3322	)	,
(	3314	)	,
(	3305	)	,
(	3297	)	,
(	3289	)	,
(	3281	)	,
(	3273	)	,
(	3265	)	,
(	3257	)	,
(	3249	)	,
(	3242	)	,
(	3234	)	,
(	3226	)	,
(	3218	)	,
(	3210	)	,
(	3203	)	,
(	3195	)	,
(	3187	)	,
(	3179	)	,
(	3172	)	,
(	3164	)	,
(	3157	)	,
(	3149	)	,
(	3142	)	,
(	3134	)	,
(	3127	)	,
(	3119	)	,
(	3112	)	,
(	3104	)	,
(	3097	)	,
(	3089	)	,
(	3082	)	,
(	3075	)	,
(	3068	)	,
(	3060	)	,
(	3053	)	,
(	3046	)	,
(	3039	)	,
(	3032	)	,
(	3024	)	,
(	3017	)	,
(	3010	)	,
(	3003	)	,
(	2996	)	,
(	2989	)	,
(	2982	)	,
(	2975	)	,
(	2968	)	,
(	2961	)	,
(	2955	)	,
(	2948	)	,
(	2941	)	,
(	2934	)	,
(	2927	)	,
(	2920	)	,
(	2914	)	,
(	2907	)	,
(	2900	)	,
(	2894	)	,
(	2887	)	,
(	2880	)	,
(	2874	)	,
(	2867	)	,
(	2861	)	,
(	2854	)	,
(	2848	)	,
(	2841	)	,
(	2835	)	,
(	2828	)	,
(	2822	)	,
(	2816	)	,
(	2809	)	,
(	2803	)	,
(	2796	)	,
(	2790	)	,
(	2784	)	,
(	2778	)	,
(	2771	)	,
(	2765	)	,
(	2759	)	,
(	2753	)	,
(	2747	)	,
(	2741	)	,
(	2735	)	,
(	2728	)	,
(	2722	)	,
(	2716	)	,
(	2710	)	,
(	2704	)	,
(	2698	)	,
(	2692	)	,
(	2687	)	,
(	2681	)	,
(	2675	)	,
(	2669	)	,
(	2663	)	,
(	2657	)	,
(	2651	)	,
(	2646	)	,
(	2640	)	,
(	2634	)	,
(	2629	)	,
(	2623	)	,
(	2617	)	,
(	2612	)	,
(	2606	)	,
(	2600	)	,
(	2595	)	,
(	2589	)	,
(	2584	)	,
(	2578	)	,
(	2573	)	,
(	2567	)	,
(	2562	)	,
(	2556	)	,
(	2551	)	,
(	2545	)	,
(	2540	)	,
(	2535	)	,
(	2529	)	,
(	2524	)	,
(	2519	)	,
(	2513	)	,
(	2508	)	,
(	2503	)	,
(	2498	)	,
(	2492	)	,
(	2487	)	,
(	2482	)	,
(	2477	)	,
(	2472	)	,
(	2467	)	,
(	2461	)	,
(	2456	)	,
(	2451	)	,
(	2446	)	,
(	2441	)	,
(	2436	)	,
(	2431	)	,
(	2426	)	,
(	2421	)	,
(	2416	)	,
(	2411	)	,
(	2407	)	,
(	2402	)	,
(	2397	)	,
(	2392	)	,
(	2387	)	,
(	2382	)	,
(	2378	)	,
(	2373	)	,
(	2368	)	,
(	2363	)	,
(	2359	)	,
(	2354	)	,
(	2349	)	,
(	2344	)	,
(	2340	)	,
(	2335	)	,
(	2331	)	,
(	2326	)	,
(	2321	)	,
(	2317	)	,
(	2312	)	,
(	2308	)	,
(	2303	)	,
(	2299	)	,
(	2294	)	,
(	2290	)	,
(	2285	)	,
(	2281	)	,
(	2277	)	,
(	2272	)	,
(	2268	)	,
(	2263	)	,
(	2259	)	,
(	2255	)	,
(	2250	)	,
(	2246	)	,
(	2242	)	,
(	2237	)	,
(	2233	)	,
(	2229	)	,
(	2225	)	,
(	2221	)	,
(	2216	)	,
(	2212	)	,
(	2208	)	,
(	2204	)	,
(	2200	)	,
(	2196	)	,
(	2192	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2167	)	,
(	2163	)	,
(	2159	)	,
(	2155	)	,
(	2151	)	,
(	2147	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2113	)	,
(	2109	)	,
(	2105	)	,
(	2101	)	,
(	2098	)	,
(	2094	)	,
(	2090	)	,
(	2086	)	,
(	2083	)	,
(	2079	)	,
(	2075	)	,
(	2072	)	,
(	2068	)	,
(	2064	)	,
(	2061	)	,
(	2057	)	,
(	2054	)	,
(	2050	)	,
(	2046	)	,
(	2043	)	,
(	2039	)	,
(	2036	)	,
(	2032	)	,
(	2029	)	,
(	2025	)	,
(	2022	)	,
(	2018	)	,
(	2015	)	,
(	2012	)	,
(	2008	)	,
(	2005	)	,
(	2001	)	,
(	1998	)	,
(	1995	)	,
(	1991	)	,
(	1988	)	,
(	1985	)	,
(	1981	)	,
(	1978	)	,
(	1975	)	,
(	1971	)	,
(	1968	)	,
(	1965	)	,
(	1962	)	,
(	1958	)	,
(	1955	)	,
(	1952	)	,
(	1949	)	,
(	1946	)	,
(	1942	)	,
(	1939	)	,
(	1936	)	,
(	1933	)	,
(	1930	)	,
(	1927	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1899	)	,
(	1896	)	,
(	1893	)	,
(	1890	)	,
(	1887	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1875	)	,
(	1872	)	,
(	1869	)	,
(	1866	)	,
(	1864	)	,
(	1861	)	,
(	1858	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1830	)	,
(	1827	)	,
(	1824	)	,
(	1821	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1800	)	,
(	1797	)	,
(	1794	)	,
(	1792	)	,
(	1789	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1779	)	,
(	1776	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1766	)	,
(	1763	)	,
(	1761	)	,
(	1758	)	,
(	1756	)	,
(	1753	)	,
(	1751	)	,
(	1748	)	,
(	1746	)	,
(	1743	)	,
(	1741	)	,
(	1738	)	,
(	1736	)	,
(	1734	)	,
(	1731	)	,
(	1729	)	,
(	1726	)	,
(	1724	)	,
(	1721	)	,
(	1719	)	,
(	1717	)	,
(	1714	)	,
(	1712	)	,
(	1710	)	,
(	1707	)	,
(	1705	)	,
(	1703	)	,
(	1700	)	,
(	1698	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1689	)	,
(	1686	)	,
(	1684	)	,
(	1682	)	,
(	1680	)	,
(	1677	)	,
(	1675	)	,
(	1673	)	,
(	1671	)	,
(	1668	)	,
(	1666	)	,
(	1664	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1653	)	,
(	1651	)	,
(	1649	)	,
(	1646	)	,
(	1644	)	,
(	1642	)	,
(	1640	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1632	)	,
(	1629	)	,
(	1627	)	,
(	1625	)	,
(	1623	)	,
(	1621	)	,
(	1619	)	,
(	1617	)	,
(	1615	)	,
(	1613	)	,
(	1611	)	,
(	1609	)	,
(	1607	)	,
(	1605	)	,
(	1603	)	,
(	1601	)	,
(	1599	)	,
(	1597	)	,
(	1595	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1581	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1563	)	,
(	1561	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1550	)	,
(	1548	)	,
(	1546	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1515	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1451	)	,
(	1449	)	,
(	1447	)	,
(	1446	)	,
(	1444	)	,
(	1443	)	,
(	1441	)	,
(	1439	)	,
(	1438	)	,
(	1436	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1430	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1422	)	,
(	1420	)	,
(	1419	)	,
(	1417	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1408	)	,
(	1406	)	,
(	1405	)	,
(	1403	)	,
(	1402	)	,
(	1400	)	,
(	1399	)	,
(	1397	)	,
(	1396	)	,
(	1394	)	,
(	1393	)	,
(	1391	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1385	)	,
(	1383	)	,
(	1382	)	,
(	1380	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1373	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1364	)	,
(	1363	)	,
(	1361	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1347	)	,
(	1345	)	,
(	1344	)	,
(	1342	)	,
(	1341	)	,
(	1339	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1334	)	,
(	1332	)	,
(	1331	)	,
(	1329	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1324	)	,
(	1322	)	,
(	1321	)	,
(	1319	)	,
(	1318	)	,
(	1317	)	,
(	1315	)	,
(	1314	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1308	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1282	)	,
(	1280	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1258	)	,
(	1257	)	,
(	1256	)	,
(	1254	)	,
(	1253	)	,
(	1252	)	,
(	1250	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1244	)	,
(	1242	)	,
(	1241	)	,
(	1240	)	,
(	1238	)	,
(	1237	)	,
(	1236	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1224	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	762	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	765	)	,
(	765	)	,
(	765	)	,
(	766	)	,
(	766	)	,
(	766	)	,
(	767	)	,
(	767	)	,
(	767	)	,
(	768	)	,
(	768	)	,
(	768	)	,
(	769	)	,
(	769	)	,
(	770	)	,
(	770	)	,
(	771	)	,
(	771	)	,
(	771	)	,
(	772	)	,
(	772	)	,
(	773	)	,
(	773	)	,
(	774	)	,
(	774	)	,
(	775	)	,
(	776	)	,
(	776	)	,
(	777	)	,
(	777	)	,
(	778	)	,
(	779	)	,
(	779	)	,
(	780	)	,
(	780	)	,
(	781	)	,
(	782	)	,
(	782	)	,
(	783	)	,
(	784	)	,
(	785	)	,
(	785	)	,
(	786	)	,
(	787	)	,
(	788	)	,
(	788	)	,
(	789	)	,
(	790	)	,
(	791	)	,
(	792	)	,
(	792	)	,
(	793	)	,
(	794	)	,
(	795	)	,
(	796	)	,
(	797	)	,
(	798	)	,
(	799	)	,
(	800	)	,
(	801	)	,
(	802	)	,
(	803	)	,
(	804	)	,
(	805	)	,
(	806	)	,
(	807	)	,
(	808	)	,
(	809	)	,
(	810	)	,
(	811	)	,
(	812	)	,
(	813	)	,
(	814	)	,
(	815	)	,
(	817	)	,
(	818	)	,
(	819	)	,
(	820	)	,
(	821	)	,
(	823	)	,
(	824	)	,
(	825	)	,
(	826	)	,
(	828	)	,
(	829	)	,
(	830	)	,
(	832	)	,
(	833	)	,
(	834	)	,
(	836	)	,
(	837	)	,
(	838	)	,
(	840	)	,
(	841	)	,
(	843	)	,
(	844	)	,
(	846	)	,
(	847	)	,
(	849	)	,
(	850	)	,
(	852	)	,
(	853	)	,
(	855	)	,
(	856	)	,
(	858	)	,
(	860	)	,
(	861	)	,
(	863	)	,
(	865	)	,
(	866	)	,
(	868	)	,
(	870	)	,
(	871	)	,
(	873	)	,
(	875	)	,
(	877	)	,
(	878	)	,
(	880	)	,
(	882	)	,
(	884	)	,
(	886	)	,
(	888	)	,
(	890	)	,
(	891	)	,
(	893	)	,
(	895	)	,
(	897	)	,
(	899	)	,
(	901	)	,
(	903	)	,
(	905	)	,
(	907	)	,
(	909	)	,
(	911	)	,
(	914	)	,
(	916	)	,
(	918	)	,
(	920	)	,
(	922	)	,
(	924	)	,
(	926	)	,
(	929	)	,
(	931	)	,
(	933	)	,
(	935	)	,
(	938	)	,
(	940	)	,
(	942	)	,
(	945	)	,
(	947	)	,
(	949	)	,
(	952	)	,
(	954	)	,
(	957	)	,
(	959	)	,
(	961	)	,
(	964	)	,
(	966	)	,
(	969	)	,
(	972	)	,
(	974	)	,
(	977	)	,
(	979	)	,
(	982	)	,
(	985	)	,
(	987	)	,
(	990	)	,
(	993	)	,
(	995	)	,
(	998	)	,
(	1001	)	,
(	1004	)	,
(	1006	)	,
(	1009	)	,
(	1012	)	,
(	1015	)	,
(	1018	)	,
(	1021	)	,
(	1023	)	,
(	1026	)	,
(	1029	)	,
(	1032	)	,
(	1035	)	,
(	1038	)	,
(	1041	)	,
(	1044	)	,
(	1047	)	,
(	1051	)	,
(	1054	)	,
(	1057	)	,
(	1060	)	,
(	1063	)	,
(	1066	)	,
(	1070	)	,
(	1073	)	,
(	1076	)	,
(	1079	)	,
(	1083	)	,
(	1086	)	,
(	1089	)	,
(	1093	)	,
(	1096	)	,
(	1099	)	,
(	1103	)	,
(	1106	)	,
(	1110	)	,
(	1113	)	,
(	1117	)	,
(	1120	)	,
(	1124	)	,
(	1127	)	,
(	1131	)	,
(	1135	)	,
(	1138	)	,
(	1142	)	,
(	1146	)	,
(	1149	)	,
(	1153	)	,
(	1157	)	,
(	1161	)	,
(	1164	)	,
(	1168	)	,
(	1172	)	,
(	1176	)	,
(	1180	)	,
(	1184	)	,
(	1188	)	,
(	1192	)	,
(	1196	)	,
(	1200	)	,
(	1204	)	,
(	1208	)	,
(	1212	)	,
(	1216	)	,
(	1220	)	,
(	1224	)	,
(	1229	)	,
(	1233	)	,
(	1237	)	,
(	1241	)	,
(	1246	)	,
(	1250	)	,
(	1254	)	,
(	1258	)	,
(	1263	)	,
(	1267	)	,
(	1272	)	,
(	1276	)	,
(	1281	)	,
(	1285	)	,
(	1290	)	,
(	1294	)	,
(	1299	)	,
(	1303	)	,
(	1308	)	,
(	1313	)	,
(	1317	)	,
(	1322	)	,
(	1327	)	,
(	1331	)	,
(	1336	)	,
(	1341	)	,
(	1346	)	,
(	1351	)	,
(	1356	)	,
(	1361	)	,
(	1365	)	,
(	1370	)	,
(	1375	)	,
(	1380	)	,
(	1385	)	,
(	1390	)	,
(	1396	)	,
(	1401	)	,
(	1406	)	,
(	1411	)	,
(	1416	)	,
(	1421	)	,
(	1427	)	,
(	1432	)	,
(	1437	)	,
(	1443	)	,
(	1448	)	,
(	1453	)	,
(	1459	)	,
(	1464	)	,
(	1470	)	,
(	1475	)	,
(	1481	)	,
(	1486	)	,
(	1492	)	,
(	1497	)	,
(	1503	)	,
(	1509	)	,
(	1514	)	,
(	1520	)	,
(	1526	)	,
(	1532	)	,
(	1537	)	,
(	1543	)	,
(	1549	)	,
(	1555	)	,
(	1561	)	,
(	1567	)	,
(	1573	)	,
(	1579	)	,
(	1585	)	,
(	1591	)	,
(	1597	)	,
(	1603	)	,
(	1609	)	,
(	1616	)	,
(	1622	)	,
(	1628	)	,
(	1634	)	,
(	1641	)	,
(	1647	)	,
(	1653	)	,
(	1660	)	,
(	1666	)	,
(	1673	)	,
(	1679	)	,
(	1686	)	,
(	1692	)	,
(	1699	)	,
(	1705	)	,
(	1712	)	,
(	1719	)	,
(	1725	)	,
(	1732	)	,
(	1739	)	,
(	1746	)	,
(	1752	)	,
(	1759	)	,
(	1766	)	,
(	1773	)	,
(	1780	)	,
(	1787	)	,
(	1794	)	,
(	1801	)	,
(	1808	)	,
(	1815	)	,
(	1822	)	,
(	1830	)	,
(	1837	)	,
(	1844	)	,
(	1851	)	,
(	1859	)	,
(	1866	)	,
(	1873	)	,
(	1881	)	,
(	1888	)	,
(	1896	)	,
(	1903	)	,
(	1911	)	,
(	1918	)	,
(	1926	)	,
(	1933	)	,
(	1941	)	,
(	1949	)	,
(	1956	)	,
(	1964	)	,
(	1972	)	,
(	1980	)	,
(	1988	)	,
(	1996	)	,
(	2004	)	,
(	2012	)	,
(	2020	)	,
(	2028	)	,
(	2036	)	,
(	2044	)	,
(	2052	)	,
(	2060	)	,
(	2068	)	,
(	2077	)	,
(	2085	)	,
(	2093	)	,
(	2101	)	,
(	2110	)	,
(	2118	)	,
(	2127	)	,
(	2135	)	,
(	2144	)	,
(	2152	)	,
(	2161	)	,
(	2170	)	,
(	2178	)	,
(	2187	)	,
(	2196	)	,
(	2204	)	,
(	2213	)	,
(	2222	)	,
(	2231	)	,
(	2240	)	,
(	2249	)	,
(	2258	)	,
(	2267	)	,
(	2276	)	,
(	2285	)	,
(	2294	)	,
(	2303	)	,
(	2313	)	,
(	2322	)	,
(	2331	)	,
(	2341	)	,
(	2350	)	,
(	2359	)	,
(	2369	)	,
(	2378	)	,
(	2388	)	,
(	2397	)	,
(	2407	)	,
(	2417	)	,
(	2426	)	,
(	2436	)	,
(	2446	)	,
(	2455	)	,
(	2465	)	,
(	2475	)	,
(	2485	)	,
(	2495	)	,
(	2505	)	,
(	2515	)	,
(	2525	)	,
(	2535	)	,
(	2545	)	,
(	2555	)	,
(	2566	)	,
(	2576	)	,
(	2586	)	,
(	2597	)	,
(	2607	)	,
(	2617	)	,
(	2628	)	,
(	2638	)	,
(	2649	)	,
(	2659	)	,
(	2670	)	,
(	2681	)	,
(	2691	)	,
(	2702	)	,
(	2713	)	,
(	2724	)	,
(	2735	)	,
(	2746	)	,
(	2756	)	,
(	2767	)	,
(	2778	)	,
(	2790	)	,
(	2801	)	,
(	2812	)	,
(	2823	)	,
(	2834	)	,
(	2846	)	,
(	2857	)	,
(	2868	)	,
(	2880	)	,
(	2891	)	,
(	2903	)	,
(	2914	)	,
(	2926	)	,
(	2937	)	,
(	2949	)	,
(	2961	)	,
(	2972	)	,
(	2984	)	,
(	2996	)	,
(	3008	)	,
(	3020	)	,
(	3032	)	,
(	3044	)	,
(	3056	)	,
(	3068	)	,
(	3080	)	,
(	3092	)	,
(	3104	)	,
(	3117	)	,
(	3129	)	,
(	3141	)	,
(	3154	)	,
(	3166	)	,
(	3179	)	,
(	3191	)	,
(	3204	)	,
(	3217	)	,
(	3229	)	,
(	3242	)	,
(	3255	)	,
(	3268	)	,
(	3280	)	,
(	3293	)	,
(	3306	)	,
(	3319	)	,
(	3332	)	,
(	3345	)	,
(	3358	)	,
(	3372	)	,
(	3385	)	,
(	3398	)	,
(	3411	)	,
(	3425	)	,
(	3438	)	,
(	3452	)	,
(	3465	)	,
(	3479	)	,
(	3492	)	,
(	3506	)	,
(	3520	)	,
(	3533	)	,
(	3547	)	,
(	3561	)	,
(	3575	)	,
(	3589	)	,
(	3603	)	,
(	3617	)	,
(	3631	)	,
(	3645	)	,
(	3659	)	,
(	3673	)	,
(	3688	)	,
(	3702	)	,
(	3716	)	,
(	3731	)	,
(	3745	)	,
(	3760	)	,
(	3774	)	,
(	3789	)	,
(	3804	)	,
(	3818	)	,
(	3833	)	,
(	3848	)	,
(	3863	)	,
(	3878	)	,
(	3893	)	,
(	3908	)	,
(	3923	)	,
(	3938	)	,
(	3953	)	,
(	3968	)	,
(	3983	)	,
(	3999	)	,
(	4014	)	,
(	4029	)	,
(	4045	)	,
(	4060	)	,
(	4076	)	,
(	4092	)	,
(	4107	)	,
(	4123	)	,
(	4139	)	,
(	4154	)	,
(	4170	)	,
(	4186	)	,
(	4202	)	,
(	4218	)	,
(	4234	)	,
(	4250	)	,
(	4267	)	,
(	4283	)	,
(	4299	)	,
(	4316	)	,
(	4332	)	,
(	4348	)	,
(	4365	)	,
(	4381	)	,
(	4398	)	,
(	4415	)	,
(	4431	)	,
(	4448	)	,
(	4465	)	,
(	4482	)	,
(	4499	)	,
(	4516	)	,
(	4533	)	,
(	4550	)	,
(	4567	)	,
(	4584	)	,
(	4602	)	,
(	4619	)	,
(	4636	)	,
(	4654	)	,
(	4671	)	,
(	4689	)	,
(	4706	)	,
(	4724	)	,
(	4742	)	,
(	4759	)	,
(	4777	)	,
(	4795	)	,
(	4813	)	,
(	4831	)	,
(	4849	)	,
(	4867	)	,
(	4885	)	,
(	4903	)	,
(	4922	)	,
(	4940	)	,
(	4958	)	,
(	4977	)	,
(	4995	)	,
(	5014	)	,
(	5032	)	,
(	5051	)	,
(	5070	)	,
(	5088	)	,
(	5107	)	,
(	5126	)	,
(	5145	)	,
(	5164	)	,
(	5183	)	,
(	5202	)	,
(	5221	)	,
(	5241	)	,
(	5260	)	,
(	5279	)	,
(	5299	)	,
(	5318	)	,
(	5338	)	,
(	5357	)	,
(	5377	)	,
(	5397	)	,
(	5416	)	,
(	5436	)	,
(	5456	)	,
(	5476	)	,
(	5496	)	,
(	5516	)	,
(	5536	)	,
(	5556	)	,
(	5577	)	,
(	5597	)	,
(	5617	)	,
(	5638	)	,
(	5658	)	,
(	5679	)	,
(	5699	)	,
(	5720	)	,
(	5741	)	,
(	5762	)	,
(	5783	)	,
(	5803	)	,
(	5824	)	,
(	5845	)	,
(	5867	)	,
(	5888	)	,
(	5909	)	,
(	5930	)	,
(	5952	)	,
(	5973	)	,
(	5994	)	,
(	6016	)	,
(	6038	)	,
(	6059	)	,
(	6081	)	,
(	6103	)	,
(	6125	)	,
(	6147	)	,
(	6169	)	,
(	6191	)	,
(	6213	)	,
(	6235	)	,
(	6257	)	,
(	6279	)	,
(	6302	)	,
(	6324	)	,
(	6347	)	,
(	6369	)	,
(	6392	)	,
(	6415	)	,
(	6437	)	,
(	6460	)	,
(	6483	)	,
(	6506	)	,
(	6529	)	,
(	6552	)	,
(	6575	)	,
(	6598	)	,
(	6622	)	,
(	6645	)	,
(	6668	)	,
(	6692	)	,
(	6715	)	,
(	6739	)	,
(	6763	)	,
(	6787	)	,
(	6810	)	,
(	6834	)	,
(	6858	)	,
(	6882	)	,
(	6906	)	,
(	6930	)	,
(	6955	)	,
(	6979	)	,
(	7003	)	,
(	7028	)	,
(	7052	)	,
(	7077	)	,
(	7101	)	,
(	7126	)	,
(	7151	)	,
(	7176	)	,
(	7200	)	,
(	7225	)	,
(	7250	)	,
(	7276	)	,
(	7301	)	,
(	7326	)	,
(	7351	)	,
(	7377	)	,
(	7402	)	,
(	7428	)	,
(	7453	)	,
(	7479	)	,
(	7505	)	,
(	7530	)	,
(	7556	)	,
(	7582	)	,
(	7608	)	,
(	7634	)	,
(	7660	)	,
(	7687	)	,
(	7713	)	,
(	7739	)	,
(	7766	)	,
(	7792	)	,
(	7819	)	,
(	7846	)	,
(	7872	)	,
(	7899	)	,
(	7926	)	,
(	7953	)	,
(	7980	)	,
(	8007	)	,
(	8034	)	,
(	8061	)	,
(	8089	)	,
(	8116	)	,
(	8144	)	,
(	8171	)	,
(	8199	)	,
(	8226	)	,
(	8254	)	,
(	8282	)	,
(	8310	)	,
(	8338	)	,
(	8366	)	,
(	8394	)	,
(	8422	)	,
(	8450	)	,
(	8479	)	,
(	8507	)	,
(	8536	)	,
(	8564	)	,
(	8593	)	,
(	8622	)	,
(	8650	)	,
(	8679	)	,
(	8708	)	,
(	8737	)	,
(	8766	)	,
(	8796	)	,
(	8825	)	,
(	8854	)	,
(	8883	)	,
(	8913	)	,
(	8943	)	,
(	8972	)	,
(	9002	)	,
(	9032	)	,
(	9062	)	,
(	9091	)	,
(	9121	)	,
(	9152	)	,
(	9182	)	,
(	9212	)	,
(	9242	)	,
(	9273	)	,
(	9303	)	,
(	9334	)	,
(	9364	)	,
(	9395	)	,
(	9426	)	,
(	9457	)	,
(	9488	)	,
(	9519	)	,
(	9550	)	,
(	9581	)	,
(	9612	)	,
(	9644	)	,
(	9675	)	,
(	9707	)	,
(	9738	)	,
(	9770	)	,
(	9802	)	,
(	9834	)	,
(	9866	)	,
(	9898	)	,
(	9930	)	,
(	9962	)	,
(	9994	)	,
(	10026	)	,
(	10059	)	,
(	10091	)	,
(	10124	)	,
(	10157	)	,
(	10189	)	,
(	10222	)	,
(	10255	)	,
(	10288	)	,
(	10321	)	,
(	10354	)	,
(	10387	)	,
(	10421	)	,
(	10454	)	,
(	10488	)	,
(	10521	)	,
(	10555	)	,
(	10589	)	,
(	10622	)	,
(	10656	)	,
(	10690	)	,
(	10724	)	,
(	10758	)	,
(	10793	)	,
(	10827	)	,
(	10861	)	,
(	10896	)	,
(	10931	)	,
(	10965	)	,
(	11000	)	,
(	11035	)	,
(	11070	)	,
(	11105	)	,
(	11140	)	,
(	11175	)	,
(	11210	)	,
(	11246	)	,
(	11281	)	,
(	11316	)	,
(	11352	)	,
(	11388	)	,
(	11424	)	,
(	11459	)	,
(	11495	)	,
(	11531	)	,
(	11568	)	,
(	11604	)	,
(	11640	)	,
(	11676	)	,
(	11713	)	,
(	11749	)	,
(	11786	)	,
(	11823	)	,
(	11860	)	,
(	11897	)	,
(	11934	)	,
(	11971	)	,
(	12008	)	,
(	12045	)	,
(	12083	)	,
(	12120	)	,
(	12158	)	,
(	12195	)	,
(	12233	)	,
(	12271	)	,
(	12309	)	,
(	12347	)	,
(	12385	)	,
(	12423	)	,
(	12461	)	,
(	12500	)	,
(	12538	)	,
(	12577	)	,
(	12615	)	,
(	12654	)	,
(	12693	)	,
(	12732	)	,
(	12771	)	,
(	12810	)	,
(	12849	)	,
(	12888	)	,
(	12928	)	,
(	12967	)	,
(	13007	)	,
(	13046	)	,
(	13086	)	,
(	13126	)	,
(	13166	)	,
(	13206	)	,
(	13246	)	,
(	13286	)	,
(	13326	)	,
(	13367	)	,
(	13407	)	,
(	13448	)	,
(	13488	)	,
(	13529	)	,
(	13570	)	,
(	13611	)	,
(	13652	)	,
(	13693	)	,
(	13735	)	,
(	13776	)	,
(	13817	)	,
(	13859	)	,
(	13900	)	,
(	13942	)	,
(	13984	)	,
(	14026	)	,
(	14068	)	,
(	14110	)	,
(	14152	)	,
(	14195	)	,
(	14237	)	,
(	14279	)	,
(	14322	)	,
(	14365	)	,
(	14408	)	,
(	14450	)	,
(	14493	)	,
(	14537	)	,
(	14580	)	,
(	14623	)	,
(	14666	)	,
(	14710	)	,
(	14753	)	,
(	14797	)	,
(	14841	)	,
(	14885	)	,
(	14929	)	,
(	14973	)	,
(	15017	)	,
(	15061	)	,
(	15106	)	,
(	15150	)	,
(	15195	)	,
(	15239	)	,
(	15284	)	,
(	15329	)	,
(	15374	)	,
(	15419	)	,
(	15464	)	,
(	15509	)	,
(	15555	)	,
(	15600	)	,
(	15646	)	,
(	15692	)	,
(	15737	)	,
(	15783	)	,
(	15829	)	,
(	15875	)	,
(	15922	)	,
(	15968	)	,
(	16014	)	,
(	16061	)	,
(	16107	)	,
(	16154	)	,
(	16201	)	,
(	16248	)	,
(	16295	)	,
(	16342	)	,
(	16389	)	,
(	16437	)	,
(	16484	)	,
(	16532	)	,
(	16579	)	,
(	16627	)	,
(	16675	)	,
(	16723	)	,
(	16771	)	,
(	16819	)	,
(	16867	)	,
(	16916	)	,
(	16964	)	,
(	17013	)	,
(	17061	)	,
(	17110	)	,
(	17159	)	,
(	17208	)	,
(	17257	)	,
(	17307	)	,
(	17356	)	,
(	17405	)	,
(	17455	)	,
(	17505	)	,
(	17554	)	,
(	17604	)	,
(	17654	)	,
(	17704	)	,
(	17755	)	,
(	17805	)	,
(	17855	)	,
(	17906	)	,
(	17956	)	,
(	18007	)	,
(	18058	)	,
(	18109	)	,
(	18160	)	,
(	18211	)	,
(	18263	)	,
(	18314	)	,
(	18365	)	,
(	18417	)	,
(	18469	)	,
(	18521	)	,
(	18573	)	,
(	18625	)	,
(	18677	)	,
(	18729	)	,
(	18782	)	,
(	18834	)	,
(	18887	)	,
(	18939	)	,
(	18992	)	,
(	19045	)	,
(	19098	)	,
(	19152	)	,
(	19205	)	,
(	19258	)	,
(	19312	)	,
(	19365	)	,
(	19419	)	,
(	19473	)	,
(	19527	)	,
(	19581	)	,
(	19635	)	,
(	19690	)	,
(	19744	)	,
(	19799	)	,
(	19853	)	,
(	19908	)	,
(	19963	)	,
(	20018	)	,
(	20073	)	,
(	20128	)	,
(	20184	)	,
(	20239	)	,
(	20295	)	,
(	20350	)	,
(	20406	)	,
(	20462	)	,
(	20518	)	,
(	20574	)	,
(	20631	)	,
(	20687	)	,
(	20744	)	,
(	20800	)	,
(	20857	)	,
(	20914	)	,
(	20971	)	,
(	21028	)	,
(	21085	)	,
(	21143	)	,
(	21200	)	,
(	21258	)	,
(	21315	)	,
(	21373	)	,
(	21431	)	,
(	21489	)	,
(	21547	)	,
(	21606	)	,
(	21664	)	,
(	21722	)	,
(	21781	)	,
(	21840	)	,
(	21899	)	,
(	21958	)	,
(	22017	)	,
(	22076	)	,
(	22136	)	,
(	22195	)	,
(	22255	)	,
(	22314	)	,
(	22374	)	,
(	22434	)	,
(	22494	)	,
(	22555	)	,
(	22615	)	,
(	22675	)	,
(	22736	)	,
(	22797	)	,
(	22858	)	,
(	22918	)	,
(	22980	)	,
(	23041	)	,
(	23102	)	,
(	23164	)	,
(	23225	)	,
(	23287	)	,
(	23349	)	,
(	23411	)	,
(	23473	)	,
(	23535	)	,
(	23597	)	,
(	23660	)	,
(	23722	)	,
(	23785	)	,
(	23848	)	,
(	23911	)	,
(	23974	)	,
(	24037	)	,
(	24100	)	,
(	24164	)	,
(	24227	)	,
(	24291	)	,
(	24355	)	,
(	24419	)	,
(	24483	)	,
(	24547	)	,
(	24611	)	,
(	24676	)	,
(	24741	)	,
(	24805	)	,
(	24870	)	,
(	24935	)	,
(	25000	)	,
(	25065	)	,
(	25131	)	,
(	25196	)	,
(	25262	)	,
(	25328	)	,
(	25394	)	,
(	25460	)	,
(	25526	)	,
(	25592	)	,
(	25658	)	,
(	25725	)	,
(	25792	)	,
(	25858	)	,
(	25925	)	,
(	25992	)	,
(	26060	)	,
(	26127	)	,
(	26194	)	,
(	26262	)	,
(	26330	)	,
(	26397	)	,
(	26465	)	,
(	26534	)	,
(	26602	)	,
(	26670	)	,
(	26739	)	,
(	26807	)	,
(	26876	)	,
(	26945	)	,
(	27014	)	,
(	27083	)	,
(	27153	)	,
(	27222	)	,
(	27292	)	,
(	27361	)	,
(	27431	)	,
(	27501	)	,
(	27571	)	,
(	27641	)	,
(	27712	)	,
(	27782	)	,
(	27853	)	,
(	27924	)	,
(	27995	)	,
(	28066	)	,
(	28137	)	,
(	28208	)	,
(	28280	)	,
(	28351	)	,
(	28423	)	,
(	28495	)	,
(	28567	)	,
(	28639	)	,
(	28712	)	,
(	28784	)	,
(	28857	)	,
(	28929	)	,
(	29002	)	,
(	29075	)	,
(	29148	)	,
(	29221	)	,
(	29295	)	,
(	29368	)	,
(	29442	)	,
(	29516	)	,
(	29590	)	,
(	29664	)	,
(	29738	)	,
(	29813	)	,
(	29887	)	,
(	29962	)	,
(	30037	)	,
(	30111	)	,
(	30187	)	,
(	30262	)	,
(	30337	)	,
(	30413	)	,
(	30488	)	,
(	30564	)	,
(	30640	)	,
(	30716	)	,
(	30792	)	,
(	30869	)	,
(	30945	)	,
(	31022	)	,
(	31099	)	,
(	31176	)	,
(	31253	)	,
(	31330	)	,
(	31407	)	,
(	31485	)	,
(	31562	)	,
(	31640	)	,
(	31718	)	,
(	31796	)	,
(	31874	)	,
(	31953	)	,
(	32031	)	,
(	32110	)	,
(	32189	)	,
(	32268	)	,
(	32347	)	,
(	32426	)	,
(	32505	)	,
(	32585	)	,
(	32665	)	,
(	32744	)	,
(	32824	)	,
(	32905	)	,
(	32985	)	,
(	33065	)	,
(	33146	)	,
(	33227	)	,
(	33307	)	,
(	33388	)	,
(	33470	)	,
(	33551	)	,
(	33632	)	,
(	33714	)	,
(	33796	)	,
(	33878	)	,
(	33960	)	,
(	34042	)	,
(	34124	)	,
(	34207	)	,
(	34289	)	,
(	34372	)	,
(	34455	)	,
(	34538	)	,
(	34622	)	,
(	34705	)	,
(	34789	)	,
(	34872	)	,
(	34956	)	,
(	35040	)	,
(	35124	)	,
(	35209	)	,
(	35293	)	,
(	35378	)	,
(	35462	)	,
(	35547	)	,
(	35632	)	,
(	35718	)	,
(	35803	)	,
(	35889	)	,
(	35974	)	,
(	36060	)	,
(	36146	)	,
(	36232	)	,
(	36319	)	,
(	36405	)	,
(	36492	)	,
(	36579	)	,
(	36666	)	,
(	36753	)	,
(	36840	)	,
(	36927	)	,
(	37015	)	,
(	37103	)	,
(	37190	)	,
(	37278	)	,
(	37367	)	,
(	37455	)	,
(	37543	)	,
(	37632	)	,
(	37721	)	,
(	37810	)	,
(	37899	)	,
(	37988	)	,
(	38078	)	,
(	38167	)	,
(	38257	)	,
(	38347	)	,
(	38437	)	,
(	38527	)	,
(	38618	)	,
(	38708	)	,
(	38799	)	,
(	38890	)	,
(	38981	)	,
(	39072	)	,
(	39164	)	,
(	39255	)	,
(	39347	)	,
(	39439	)	,
(	39531	)	,
(	39623	)	,
(	39715	)	,
(	39808	)	,
(	39900	)	,
(	39993	)	,
(	40086	)	,
(	40179	)	,
(	40272	)	,
(	40366	)	,
(	40460	)	,
(	40553	)	,
(	40647	)	,
(	40741	)	,
(	40836	)	,
(	40930	)	,
(	41025	)	,
(	41119	)	,
(	41214	)	,
(	41309	)	,
(	41405	)	,
(	41500	)	,
(	41596	)	,
(	41692	)	,
(	41787	)	,
(	41884	)	,
(	41980	)	,
(	42076	)	,
(	42173	)	,
(	42270	)	,
(	42367	)	,
(	42464	)	,
(	42561	)	,
(	42658	)	,
(	42756	)	,
(	42854	)	,
(	42952	)	,
(	43050	)	,
(	43148	)	,
(	43246	)	,
(	43345	)	,
(	43444	)	,
(	43543	)	,
(	43642	)	,
(	43741	)	,
(	43841	)	,
(	43940	)	,
(	44040	)	,
(	44140	)	,
(	44240	)	,
(	44340	)	,
(	44441	)	,
(	44542	)	,
(	44642	)	,
(	44743	)	,
(	44844	)	,
(	44946	)	,
(	45047	)	,
(	45149	)	,
(	45251	)	,
(	45353	)	,
(	45455	)	,
(	45557	)	,
(	45660	)	,
(	45763	)	,
(	45866	)	,
(	45969	)	,
(	46072	)	,
(	46175	)	,
(	46279	)	,
(	46383	)	,
(	46487	)	,
(	46591	)	,
(	46695	)	,
(	46799	)	,
(	46904	)	,
(	47009	)	,
(	47114	)	,
(	47219	)	,
(	47324	)	,
(	47430	)	,
(	47536	)	,
(	47641	)	,
(	47747	)	,
(	47854	)	,
(	47960	)	,
(	48067	)	,
(	48173	)	,
(	48280	)	,
(	48387	)	,
(	48495	)	,
(	48602	)	,
(	48710	)	,
(	48818	)	,
(	48926	)	,
(	49034	)	,
(	49142	)	,
(	49251	)	,
(	49359	)	,
(	49468	)	,
(	49577	)	,
(	49687	)	,
(	49796	)	,
(	49906	)	,
(	50016	)	,
(	50126	)	,
(	50236	)	,
(	50346	)	,
(	50457	)	,
(	50567	)	,
(	50678	)	,
(	50789	)	,
(	50901	)	,
(	51012	)	,
(	51124	)	,
(	51235	)	,
(	51347	)	,
(	51460	)	,
(	51572	)	,
(	51685	)	,
(	51797	)	,
(	51910	)	,
(	52023	)	,
(	52137	)	,
(	52250	)	,
(	52364	)	,
(	52478	)	,
(	52592	)	,
(	52706	)	,
(	52820	)	,
(	52935	)	,
(	53050	)	,
(	53165	)	,
(	53280	)	,
(	53395	)	,
(	53511	)	,
(	53626	)	,
(	53742	)	,
(	53858	)	,
(	53975	)	,
(	54091	)	,
(	54208	)	,
(	54324	)	,
(	54441	)	,
(	54559	)	,
(	54676	)	,
(	54794	)	,
(	54911	)	,
(	55029	)	,
(	55148	)	,
(	55266	)	,
(	55385	)	,
(	55503	)	,
(	55622	)	,
(	55741	)	,
(	55861	)	,
(	55980	)	,
(	56100	)	,
(	56220	)	,
(	56340	)	,
(	56460	)	,
(	56581	)	,
(	56701	)	,
(	56822	)	,
(	56943	)	,
(	57064	)	,
(	57186	)	,
(	57307	)	,
(	57429	)	,
(	57551	)	,
(	57673	)	,
(	57796	)	,
(	57918	)	,
(	58041	)	,
(	58164	)	,
(	58287	)	,
(	58411	)	,
(	58534	)	,
(	58658	)	,
(	58782	)	,
(	58906	)	,
(	59031	)	,
(	59155	)	,
(	59280	)	,
(	59405	)	,
(	59530	)	,
(	59655	)	,
(	59781	)	,
(	59907	)	,
(	60033	)	,
(	60159	)	,
(	60285	)	,
(	60412	)	,
(	60538	)	,
(	60665	)	,
(	60792	)	,
(	60920	)	,
(	61047	)	,
(	61175	)	,
(	61303	)	,
(	61431	)	,
(	61559	)	,
(	61688	)	,
(	61817	)	,
(	61946	)	,
(	62075	)	,
(	62204	)	,
(	62334	)	,
(	62463	)	,
(	62593	)	,
(	62724	)	,
(	62854	)	,
(	62984	)	,
(	63115	)	,
(	63246	)	,
(	63377	)	,
(	63509	)	,
(	63640	)	,
(	63772	)	,
(	63904	)	,
(	64036	)	,
(	64169	)	,
(	64301	)	,
(	64434	)	,
(	64567	)	,
(	64700	)	,
(	64834	)	,
(	64967	)	,
(	65101	)	,
(	65235	)	,
(	65370	)	,
(	65504	)	,
(	65639	)	,
(	65774	)	,
(	65909	)	,
(	66044	)	,
(	66179	)	,
(	66315	)	,
(	66451	)	,
(	66587	)	,
(	66724	)	,
(	66860	)	,
(	66997	)	,
(	67134	)	,
(	67271	)	,
(	67408	)	,
(	67546	)	,
(	67684	)	,
(	67822	)	,
(	67960	)	,
(	68098	)	,
(	68237	)	,
(	68376	)	,
(	68515	)	,
(	68654	)	,
(	68794	)	,
(	68933	)	,
(	69073	)	,
(	69214	)	,
(	69354	)	,
(	69494	)	,
(	69635	)	,
(	69776	)	,
(	69917	)	,
(	70059	)	,
(	70200	)	,
(	70342	)	,
(	70484	)	,
(	70627	)	,
(	70769	)	,
(	70912	)	,
(	71055	)	,
(	71198	)	,
(	71341	)	,
(	71485	)	,
(	71629	)	,
(	71773	)	,
(	71917	)	,
(	72061	)	,
(	72206	)	,
(	72351	)	,
(	72496	)	,
(	72641	)	,
(	72787	)	,
(	72932	)	,
(	73078	)	,
(	73225	)	,
(	73371	)	,
(	73518	)	,
(	73665	)	,
(	73812	)	,
(	73959	)	,
(	74106	)	,
(	74254	)	,
(	74402	)	,
(	74550	)	,
(	74699	)	,
(	74847	)	,
(	74996	)	,
(	75145	)	,
(	75294	)	,
(	75444	)	,
(	75594	)	,
(	75743	)	,
(	75894	)	,
(	76044	)	,
(	76195	)	,
(	76345	)	,
(	76497	)	,
(	76648	)	,
(	76799	)	,
(	76951	)	,
(	77103	)	,
(	77255	)	,
(	77408	)	,
(	77560	)	,
(	77713	)	,
(	77866	)	,
(	78019	)	,
(	78173	)	,
(	78327	)	,
(	78481	)	,
(	78635	)	,
(	78789	)	,
(	78944	)	,
(	79099	)	,
(	79254	)	,
(	79409	)	,
(	79565	)	,
(	79721	)	,
(	79877	)	,
(	80033	)	,
(	80190	)	,
(	80346	)	,
(	80503	)	,
(	80660	)	,
(	80818	)	,
(	80975	)	,
(	81133	)	,
(	81291	)	,
(	81450	)	,
(	81608	)	,
(	81767	)	,
(	81926	)	,
(	82085	)	,
(	82245	)	,
(	82405	)	,
(	82565	)	,
(	82725	)	,
(	82885	)	,
(	83046	)	,
(	83207	)	,
(	83368	)	,
(	83529	)	,
(	83691	)	,
(	83853	)	,
(	84015	)	,
(	84177	)	,
(	84339	)	,
(	84502	)	,
(	84665	)	,
(	84828	)	,
(	84992	)	,
(	85156	)	,
(	85320	)	,
(	85484	)	,
(	85648	)	,
(	85813	)	,
(	85978	)	,
(	86143	)	,
(	86308	)	,
(	86474	)	,
(	86640	)	,
(	86806	)	,
(	86972	)	,
(	87139	)	,
(	87305	)	,
(	87472	)	,
(	87640	)	,
(	87807	)	,
(	87975	)	,
(	88143	)	,
(	88311	)	,
(	88480	)	,
(	88648	)	,
(	88817	)	,
(	88986	)	,
(	89156	)	,
(	89326	)	,
(	89496	)	,
(	89666	)	,
(	89836	)	,
(	90007	)	,
(	90178	)	,
(	90349	)	,
(	90520	)	,
(	90692	)	,
(	90864	)	,
(	91036	)	,
(	91208	)	,
(	91381	)	,
(	91554	)	,
(	91727	)	,
(	91900	)	,
(	92073	)	,
(	92247	)	,
(	92421	)	,
(	92596	)	,
(	92770	)	,
(	92945	)	,
(	93120	)	,
(	93295	)	,
(	93471	)	,
(	93647	)	,
(	93823	)	,
(	93999	)	,
(	94176	)	,
(	94352	)	,
(	94529	)	,
(	94707	)	,
(	94884	)	,
(	95062	)	,
(	95240	)	,
(	95418	)	,
(	95597	)	,
(	95776	)	,
(	95955	)	,
(	96134	)	,
(	96314	)	,
(	96493	)	,
(	96673	)	,
(	96854	)	,
(	97034	)	,
(	97215	)	,
(	97396	)	,
(	97577	)	,
(	97759	)	,
(	97941	)	,
(	98123	)	,
(	98305	)	,
(	98488	)	,
(	98670	)	,
(	98853	)	,
(	99037	)	,
(	99220	)	,
(	99404	)	,
(	99588	)	,
(	99773	)	,
(	99957	)	,
(	100142	)	,
(	100327	)	,
(	100513	)	,
(	100698	)	,
(	100884	)	,
(	101070	)	,
(	101257	)	,
(	101443	)	,
(	101630	)	,
(	101817	)	,
(	102005	)	,
(	102192	)	,
(	102380	)	,
(	102569	)	,
(	102757	)	,
(	102946	)	,
(	103135	)	,
(	103324	)	,
(	103514	)	,
(	103703	)	,
(	103893	)	,
(	104084	)	,
(	104274	)	,
(	104465	)	,
(	104656	)	,
(	104847	)	,
(	105039	)	,
(	105231	)	,
(	105423	)	,
(	105615	)	,
(	105808	)	,
(	106001	)	,
(	106194	)	,
(	106387	)	,
(	106581	)	,
(	106775	)	,
(	106969	)	,
(	107164	)	,
(	107359	)	,
(	107554	)	,
(	107749	)	,
(	107944	)	,
(	108140	)	,
(	108336	)	,
(	108533	)	,
(	108729	)	,
(	108926	)	,
(	109123	)	,
(	109321	)	,
(	109518	)	,
(	109716	)	,
(	109915	)	,
(	110113	)	,
(	110312	)	,
(	110511	)	,
(	110710	)	,
(	110910	)	,
(	111109	)	,
(	111310	)	,
(	111510	)	,
(	111711	)	,
(	111911	)	,
(	112113	)	,
(	112314	)	,
(	112516	)	,
(	112718	)	,
(	112920	)	,
(	113123	)	,
(	113325	)	,
(	113528	)	,
(	113732	)	,
(	113935	)	,
(	114139	)	,
(	114344	)	,
(	114548	)	,
(	114753	)	,
(	114958	)	,
(	115163	)	,
(	115369	)	,
(	115574	)	,
(	115780	)	,
(	115987	)	,
(	116193	)	,
(	116400	)	,
(	116608	)	,
(	116815	)	,
(	117023	)	,
(	117231	)	,
(	117439	)	,
(	117648	)	,
(	117857	)	,
(	118066	)	,
(	118275	)	,
(	118485	)	,
(	118695	)	,
(	118905	)	,
(	119115	)	,
(	119326	)	,
(	119537	)	,
(	119749	)	,
(	119960	)	,
(	120172	)	,
(	120385	)	,
(	120597	)	,
(	120810	)	,
(	121023	)	,
(	121236	)	,
(	121450	)	,
(	121664	)	,
(	121878	)	,
(	122092	)	,
(	122307	)	,
(	122522	)	,
(	122737	)	,
(	122953	)	,
(	123169	)	,
(	123385	)	,
(	123601	)	,
(	123818	)	,
(	124035	)	,
(	124252	)	,
(	124470	)	,
(	124688	)	,
(	124906	)	,
(	125124	)	,
(	125343	)	,
(	125562	)	,
(	125781	)	,
(	126001	)	,
(	126221	)	,
(	126441	)	,
(	126661	)	,
(	126882	)	,
(	127103	)	,
(	127324	)	,
(	127546	)	,
(	127768	)	,
(	127990	)	,
(	128213	)	,
(	128435	)	,
(	128658	)	,
(	128882	)	,
(	129105	)	,
(	129329	)	,
(	129553	)	,
(	129778	)	,
(	130003	)	,
(	130228	)	,
(	130453	)	,
(	130679	)	,
(	130905	)	,
(	131131	)	,
(	131358	)	,
(	131584	)	,
(	131812	)	,
(	132039	)	,
(	132267	)	,
(	132495	)	,
(	132723	)	,
(	132952	)	,
(	133180	)	,
(	133410	)	,
(	133639	)	,
(	133869	)	,
(	134099	)	,
(	134329	)	,
(	134560	)	,
(	134791	)	,
(	135022	)	,
(	135254	)	,
(	135486	)	,
(	135718	)	,
(	135950	)	,
(	136183	)	,
(	136416	)	,
(	136649	)	,
(	136883	)	,
(	137117	)	,
(	137351	)	,
(	137586	)	,
(	137820	)	,
(	138056	)	,
(	138291	)	,
(	138527	)	,
(	138763	)	,
(	138999	)	,
(	139236	)	,
(	139473	)	,
(	139710	)	,
(	139948	)	,
(	140185	)	,
(	140424	)	,
(	140662	)	,
(	140901	)	,
(	141140	)	,
(	141379	)	,
(	141619	)	,
(	141859	)	,
(	142099	)	,
(	142340	)	,
(	142581	)	,
(	142822	)	,
(	143063	)	,
(	143305	)	,
(	143547	)	,
(	143790	)	,
(	144032	)	,
(	144275	)	,
(	144519	)	,
(	144762	)	,
(	145006	)	,
(	145250	)	,
(	145495	)	,
(	145740	)	,
(	145985	)	,
(	146231	)	,
(	146476	)	,
(	146723	)	,
(	146969	)	,
(	147216	)	,
(	147463	)	,
(	147710	)	,
(	147958	)	,
(	148206	)	,
(	148454	)	,
(	148703	)	,
(	148951	)	,
(	149201	)	,
(	149450	)	,
(	149700	)	,
(	149950	)	,
(	150201	)	,
(	150451	)	,
(	150703	)	,
(	150954	)	,
(	151206	)	,
(	151458	)	,
(	151710	)	,
(	151963	)	,
(	152216	)	,
(	152469	)	,
(	152723	)	,
(	152977	)	,
(	153231	)	,
(	153485	)	,
(	153740	)	,
(	153995	)	,
(	154251	)	,
(	154507	)	,
(	154763	)	,
(	155019	)	,
(	155276	)	,
(	155533	)	,
(	155791	)	,
(	156048	)	,
(	156307	)	,
(	156565	)	,
(	156824	)	,
(	157083	)	,
(	157342	)	,
(	157602	)	,
(	157862	)	,
(	158122	)	,
(	158383	)	,
(	158643	)	,
(	158905	)	,
(	159166	)	,
(	159428	)	,
(	159690	)	,
(	159953	)	,
(	160216	)	,
(	160479	)	,
(	160743	)	,
(	161006	)	,
(	161271	)	,
(	161535	)	,
(	161800	)	,
(	162065	)	,
(	162331	)	,
(	162596	)	,
(	162863	)	,
(	163129	)	,
(	163396	)	,
(	163663	)	,
(	163930	)	,
(	164198	)	,
(	164466	)	,
(	164735	)	,
(	165003	)	,
(	165272	)	,
(	165542	)	,
(	165811	)	,
(	166082	)	,
(	166352	)	,
(	166623	)	,
(	166894	)	,
(	167165	)	,
(	167437	)	,
(	167709	)	,
(	167981	)	,
(	168254	)	,
(	168527	)	,
(	168800	)	,
(	169074	)	,
(	169348	)	,
(	169622	)	,
(	169897	)	,
(	170172	)	,
(	170447	)	,
(	170723	)	,
(	170999	)	,
(	171275	)	,
(	171552	)	,
(	171829	)	,
(	172107	)	,
(	172384	)	,
(	172662	)	,
(	172941	)	,
(	173219	)	,
(	173498	)	,
(	173778	)	,
(	174057	)	,
(	174338	)	,
(	174618	)	,
(	174899	)	,
(	175180	)	,
(	175461	)	,
(	175743	)	,
(	176025	)	,
(	176307	)	,
(	176590	)	,
(	176873	)	,
(	177157	)	,
(	177440	)	,
(	177725	)	,
(	178009	)	,
(	178294	)	,
(	178579	)	,
(	178864	)	,
(	179150	)	,
(	179436	)	,
(	179723	)	,
(	180010	)	,
(	180297	)	,
(	180585	)	,
(	180872	)	,
(	181161	)	,
(	181449	)	,
(	181738	)	,
(	182027	)	,
(	182317	)	,
(	182607	)	,
(	182897	)	,
(	183188	)	,
(	183479	)	,
(	183770	)	,
(	184062	)	,
(	184354	)	,
(	184646	)	,
(	184939	)	,
(	185232	)	,
(	185525	)	,
(	185819	)	,
(	186113	)	,
(	186408	)	,
(	186702	)	,
(	186998	)	,
(	187293	)	,
(	187589	)	,
(	187885	)	,
(	188182	)	,
(	188479	)	,
(	188776	)	,
(	189073	)	,
(	189371	)	,
(	189670	)	,
(	189968	)	,
(	190267	)	,
(	190567	)	,
(	190866	)	,
(	191167	)	,
(	191467	)	,
(	191768	)	,
(	192069	)	,
(	192370	)	,
(	192672	)	,
(	192974	)	,
(	193277	)	,
(	193580	)	,
(	193883	)	,
(	194187	)	,
(	194491	)	,
(	194795	)	,
(	195100	)	,
(	195405	)	,
(	195710	)	,
(	196016	)	,
(	196322	)	,
(	196628	)	,
(	196935	)	,
(	197242	)	,
(	197550	)	,
(	197858	)	,
(	198166	)	,
(	198475	)	,
(	198784	)	,
(	199093	)	,
(	199403	)	,
(	199713	)	,
(	200023	)	,
(	200334	)	,
(	200645	)	,
(	200957	)	,
(	201269	)	,
(	201581	)	,
(	201893	)	,
(	202206	)	,
(	202520	)	,
(	202833	)	,
(	203147	)	,
(	203462	)	,
(	203777	)	,
(	204092	)	,
(	204407	)	,
(	204723	)	,
(	205039	)	,
(	205356	)	,
(	205673	)	,
(	205990	)	,
(	206308	)	,
(	206626	)	,
(	206944	)	,
(	207263	)	,
(	207582	)	,
(	207902	)	,
(	208222	)	,
(	208542	)	,
(	208863	)	,
(	209184	)	,
(	209505	)	,
(	209827	)	,
(	210149	)	,
(	210472	)	,
(	210794	)	,
(	211118	)	,
(	211441	)	,
(	211765	)	,
(	212090	)	,
(	212414	)	,
(	212739	)	,
(	213065	)	,
(	213391	)	,
(	213717	)	,
(	214043	)	,
(	214370	)	,
(	214698	)	,
(	215025	)	,
(	215354	)	,
(	215682	)	,
(	216011	)	,
(	216340	)	,
(	216670	)	,
(	217000	)	,
(	217330	)	,
(	217661	)	,
(	217992	)	,
(	218323	)	,
(	218655	)	,
(	218987	)	,
(	219320	)	,
(	219653	)	,
(	219986	)	,
(	220320	)	,
(	220654	)	,
(	220988	)	,
(	221323	)	,
(	221659	)	,
(	221994	)	,
(	222330	)	,
(	222667	)	,
(	223003	)	,
(	223340	)	,
(	223678	)	,
(	224016	)	,
(	224354	)	,
(	224693	)	,
(	225032	)	,
(	225371	)	,
(	225711	)	,
(	226051	)	,
(	226392	)	,
(	226733	)	,
(	227074	)	,
(	227416	)	,
(	227758	)	,
(	228101	)	,
(	228444	)	,
(	228787	)	,
(	229131	)	,
(	229475	)	,
(	229819	)	,
(	230164	)	,
(	230509	)	,
(	230855	)	,
(	231201	)	,
(	231547	)	,
(	231894	)	,
(	232241	)	,
(	232589	)	,
(	232937	)	,
(	233285	)	,
(	233634	)	,
(	233983	)	,
(	234332	)	,
(	234682	)	,
(	235033	)	,
(	235383	)	,
(	235734	)	,
(	236086	)	,
(	236438	)	,
(	236790	)	,
(	237143	)	,
(	237496	)	,
(	237849	)	,
(	238203	)	,
(	238557	)	,
(	238912	)	,
(	239267	)	,
(	239622	)	,
(	239978	)	,
(	240334	)	,
(	240691	)	,
(	241048	)	,
(	241405	)	,
(	241763	)	,
(	242121	)	,
(	242480	)	,
(	242839	)	,
(	243198	)	,
(	243558	)	,
(	243918	)	,
(	244278	)	,
(	244639	)	,
(	245001	)	,
(	245362	)	,
(	245725	)	,
(	246087	)	,
(	246450	)	,
(	246813	)	,
(	247177	)	,
(	247541	)	,
(	247906	)	,
(	248271	)	,
(	248636	)	,
(	249002	)	,
(	249368	)	,
(	249735	)	,
(	250102	)	,
(	250469	)	,
(	250837	)	,
(	251205	)	,
(	251574	)	,
(	251943	)	,
(	252312	)	,
(	252682	)	,
(	253052	)	,
(	253423	)	,
(	253794	)	,
(	254165	)	,
(	254537	)	,
(	254909	)	,
(	255282	)	,
(	255655	)	,
(	256029	)	,
(	256403	)	,
(	256777	)	,
(	257152	)	,
(	257527	)	,
(	257902	)	,
(	258278	)	,
(	258654	)	,
(	259031	)	,
(	259408	)	,
(	259786	)	,
(	260164	)	,
(	260542	)	,
(	260921	)	,
(	261300	)	,
(	261680	)	,
(	262060	)	,
(	262440	)	,
(	262821	)	,
(	263203	)	,
(	263584	)	,
(	263966	)	,
(	264349	)	,
(	264732	)	,
(	265115	)	,
(	265499	)	,
(	265883	)	,
(	266268	)	,
(	266653	)	,
(	267038	)	,
(	267424	)	,
(	267811	)	,
(	268197	)	,
(	268584	)	,
(	268972	)	,
(	269360	)	,
(	269748	)	,
(	270137	)	,
(	270526	)	,
(	270916	)	,
(	271306	)	,
(	271696	)	,
(	272087	)	,
(	272479	)	,
(	272870	)	,
(	273262	)	,
(	273655	)	,
(	274048	)	,
(	274441	)	,
(	274835	)	,
(	275230	)	,
(	275624	)	,
(	276019	)	,
(	276415	)	,
(	276811	)	,
(	277207	)	,
(	277604	)	,
(	278001	)	,
(	278399	)	,
(	278797	)	,
(	279196	)	,
(	279594	)	,
(	279994	)	,
(	280394	)	,
(	280794	)	,
(	281195	)	,
(	281596	)	,
(	281997	)	,
(	282399	)	,
(	282801	)	,
(	283204	)	,
(	283607	)	,
(	284011	)	,
(	284415	)	,
(	284820	)	,
(	285225	)	,
(	285630	)	,
(	286036	)	,
(	286442	)	,
(	286849	)	,
(	287256	)	,
(	287663	)	,
(	288071	)	,
(	288480	)	,
(	288889	)	,
(	289298	)	,
(	289708	)	,
(	290118	)	,
(	290528	)	,
(	290939	)	,
(	291351	)	,
(	291763	)	,
(	292175	)	,
(	292588	)	,
(	293001	)	,
(	293414	)	,
(	293829	)	,
(	294243	)	,
(	294658	)	,
(	295073	)	,
(	295489	)	,
(	295905	)	,
(	296322	)	,
(	296739	)	,
(	297157	)	,
(	297575	)	,
(	297993	)	,
(	298412	)	,
(	298832	)	,
(	299251	)	,
(	299672	)	,
(	300092	)	,
(	300513	)	,
(	300935	)	,
(	301357	)	,
(	301779	)	,
(	302202	)	,
(	302625	)	,
(	303049	)	,
(	303473	)	,
(	303898	)	,
(	304323	)	,
(	304749	)	,
(	305175	)	,
(	305601	)	,
(	306028	)	,
(	306455	)	,
(	306883	)	,
(	307311	)	,
(	307740	)	,
(	308169	)	,
(	308599	)	,
(	309029	)	,
(	309459	)	,
(	309890	)	,
(	310321	)	,
(	310753	)	,
(	311185	)	,
(	311618	)	,
(	312051	)	,
(	312485	)	,
(	312919	)	,
(	313353	)	,
(	313788	)	,
(	314224	)	,
(	314660	)	,
(	315096	)	,
(	315533	)	,
(	315970	)	,
(	316408	)	,
(	316846	)	,
(	317284	)	,
(	317723	)	,
(	318163	)	,
(	318603	)	,
(	319043	)	,
(	319484	)	,
(	319925	)	,
(	320367	)	,
(	320809	)	,
(	321252	)	,
(	321695	)	,
(	322139	)	,
(	322583	)	,
(	323027	)	,
(	323472	)	,
(	323918	)	,
(	324364	)	,
(	324810	)	,
(	325257	)	,
(	325704	)	,
(	326152	)	,
(	326600	)	,
(	327049	)	,
(	327498	)	,
(	327947	)	,
(	328397	)	,
(	328848	)	,
(	329299	)	,
(	329750	)	,
(	330202	)	,
(	330655	)	,
(	331107	)	,
(	331561	)	,
(	332015	)	,
(	332469	)	,
(	332923	)	,
(	333379	)	,
(	333834	)	,
(	334290	)	,
(	334747	)	,
(	335204	)	,
(	335661	)	,
(	336119	)	,
(	336578	)	,
(	337037	)	,
(	337496	)	,
(	337956	)	,
(	338416	)	,
(	338877	)	,
(	339338	)	,
(	339800	)	,
(	340262	)	,
(	340725	)	,
(	341188	)	,
(	341651	)	,
(	342115	)	,
(	342580	)	,
(	343045	)	,
(	343510	)	,
(	343976	)	,
(	344443	)	,
(	344910	)	,
(	345377	)	,
(	345845	)	,
(	346313	)	,
(	346782	)	,
(	347251	)	,
(	347721	)	,
(	348191	)	,
(	348662	)	,
(	349133	)	,
(	349605	)	,
(	350077	)	,
(	350549	)	,
(	351022	)	,
(	351496	)	,
(	351970	)	,
(	352444	)	,
(	352919	)	,
(	353395	)	,
(	353871	)	,
(	354347	)	,
(	354824	)	,
(	355302	)	,
(	355779	)	,
(	356258	)	,
(	356737	)	,
(	357216	)	,
(	357696	)	,
(	358176	)	,
(	358657	)	,
(	359138	)	,
(	359620	)	,
(	360102	)	,
(	360585	)	,
(	361068	)	,
(	361552	)	,
(	362036	)	,
(	362520	)	,
(	363006	)	,
(	363491	)	,
(	363977	)	,
(	364464	)	,
(	364951	)	,
(	365438	)	,
(	365926	)	,
(	366415	)	,
(	366904	)	,
(	367394	)	,
(	367884	)	,
(	368374	)	,
(	368865	)	,
(	369356	)	,
(	369848	)	,
(	370341	)	,
(	370834	)	,
(	371327	)	,
(	371821	)	,
(	372316	)	,
(	372811	)	,
(	373306	)	,
(	373802	)	,
(	374298	)	,
(	374795	)	,
(	375292	)	,
(	375790	)	,
(	376289	)	,
(	376788	)	,
(	377287	)	,
(	377787	)	,
(	378287	)	,
(	378788	)	,
(	379289	)	,
(	379791	)	,
(	380293	)	,
(	380796	)	,
(	381300	)	,
(	381803	)	,
(	382308	)	,
(	382813	)	,
(	383318	)	,
(	383824	)	,
(	384330	)	,
(	384837	)	,
(	385344	)	,
(	385852	)	,
(	386360	)	,
(	386869	)	,
(	387379	)	,
(	387888	)	,
(	388399	)	,
(	388910	)	,
);


end package LUT_pkg;
