library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4879	)	,
(	4872	)	,
(	4865	)	,
(	4858	)	,
(	4851	)	,
(	4845	)	,
(	4838	)	,
(	4831	)	,
(	4824	)	,
(	4818	)	,
(	4811	)	,
(	4804	)	,
(	4798	)	,
(	4791	)	,
(	4784	)	,
(	4777	)	,
(	4771	)	,
(	4764	)	,
(	4757	)	,
(	4751	)	,
(	4744	)	,
(	4737	)	,
(	4731	)	,
(	4724	)	,
(	4718	)	,
(	4711	)	,
(	4704	)	,
(	4698	)	,
(	4691	)	,
(	4685	)	,
(	4678	)	,
(	4671	)	,
(	4665	)	,
(	4658	)	,
(	4652	)	,
(	4645	)	,
(	4639	)	,
(	4632	)	,
(	4626	)	,
(	4619	)	,
(	4613	)	,
(	4606	)	,
(	4600	)	,
(	4593	)	,
(	4587	)	,
(	4580	)	,
(	4574	)	,
(	4567	)	,
(	4561	)	,
(	4554	)	,
(	4548	)	,
(	4542	)	,
(	4535	)	,
(	4529	)	,
(	4522	)	,
(	4516	)	,
(	4509	)	,
(	4503	)	,
(	4497	)	,
(	4490	)	,
(	4484	)	,
(	4478	)	,
(	4471	)	,
(	4465	)	,
(	4459	)	,
(	4452	)	,
(	4446	)	,
(	4440	)	,
(	4433	)	,
(	4427	)	,
(	4421	)	,
(	4414	)	,
(	4408	)	,
(	4402	)	,
(	4396	)	,
(	4389	)	,
(	4383	)	,
(	4377	)	,
(	4371	)	,
(	4364	)	,
(	4358	)	,
(	4352	)	,
(	4346	)	,
(	4340	)	,
(	4333	)	,
(	4327	)	,
(	4321	)	,
(	4315	)	,
(	4309	)	,
(	4303	)	,
(	4296	)	,
(	4290	)	,
(	4284	)	,
(	4278	)	,
(	4272	)	,
(	4266	)	,
(	4260	)	,
(	4254	)	,
(	4248	)	,
(	4241	)	,
(	4235	)	,
(	4229	)	,
(	4223	)	,
(	4217	)	,
(	4211	)	,
(	4205	)	,
(	4199	)	,
(	4193	)	,
(	4187	)	,
(	4181	)	,
(	4175	)	,
(	4169	)	,
(	4163	)	,
(	4157	)	,
(	4151	)	,
(	4145	)	,
(	4139	)	,
(	4133	)	,
(	4127	)	,
(	4121	)	,
(	4115	)	,
(	4109	)	,
(	4103	)	,
(	4097	)	,
(	4092	)	,
(	4086	)	,
(	4080	)	,
(	4074	)	,
(	4068	)	,
(	4062	)	,
(	4056	)	,
(	4050	)	,
(	4044	)	,
(	4039	)	,
(	4033	)	,
(	4027	)	,
(	4021	)	,
(	4015	)	,
(	4009	)	,
(	4004	)	,
(	3998	)	,
(	3992	)	,
(	3986	)	,
(	3980	)	,
(	3975	)	,
(	3969	)	,
(	3963	)	,
(	3957	)	,
(	3952	)	,
(	3946	)	,
(	3940	)	,
(	3934	)	,
(	3929	)	,
(	3923	)	,
(	3917	)	,
(	3912	)	,
(	3906	)	,
(	3900	)	,
(	3895	)	,
(	3889	)	,
(	3883	)	,
(	3878	)	,
(	3872	)	,
(	3866	)	,
(	3861	)	,
(	3855	)	,
(	3849	)	,
(	3844	)	,
(	3838	)	,
(	3832	)	,
(	3827	)	,
(	3821	)	,
(	3816	)	,
(	3810	)	,
(	3805	)	,
(	3799	)	,
(	3793	)	,
(	3788	)	,
(	3782	)	,
(	3777	)	,
(	3771	)	,
(	3766	)	,
(	3760	)	,
(	3755	)	,
(	3749	)	,
(	3744	)	,
(	3738	)	,
(	3733	)	,
(	3727	)	,
(	3722	)	,
(	3716	)	,
(	3711	)	,
(	3705	)	,
(	3700	)	,
(	3694	)	,
(	3689	)	,
(	3684	)	,
(	3678	)	,
(	3673	)	,
(	3667	)	,
(	3662	)	,
(	3657	)	,
(	3651	)	,
(	3646	)	,
(	3640	)	,
(	3635	)	,
(	3630	)	,
(	3624	)	,
(	3619	)	,
(	3614	)	,
(	3608	)	,
(	3603	)	,
(	3598	)	,
(	3592	)	,
(	3587	)	,
(	3582	)	,
(	3576	)	,
(	3571	)	,
(	3566	)	,
(	3560	)	,
(	3555	)	,
(	3550	)	,
(	3545	)	,
(	3539	)	,
(	3534	)	,
(	3529	)	,
(	3524	)	,
(	3518	)	,
(	3513	)	,
(	3508	)	,
(	3503	)	,
(	3498	)	,
(	3492	)	,
(	3487	)	,
(	3482	)	,
(	3477	)	,
(	3472	)	,
(	3467	)	,
(	3461	)	,
(	3456	)	,
(	3451	)	,
(	3446	)	,
(	3441	)	,
(	3436	)	,
(	3431	)	,
(	3425	)	,
(	3420	)	,
(	3415	)	,
(	3410	)	,
(	3405	)	,
(	3400	)	,
(	3395	)	,
(	3390	)	,
(	3385	)	,
(	3380	)	,
(	3375	)	,
(	3370	)	,
(	3365	)	,
(	3360	)	,
(	3355	)	,
(	3349	)	,
(	3344	)	,
(	3339	)	,
(	3334	)	,
(	3329	)	,
(	3324	)	,
(	3320	)	,
(	3315	)	,
(	3310	)	,
(	3305	)	,
(	3300	)	,
(	3295	)	,
(	3290	)	,
(	3285	)	,
(	3280	)	,
(	3275	)	,
(	3270	)	,
(	3265	)	,
(	3260	)	,
(	3255	)	,
(	3250	)	,
(	3246	)	,
(	3241	)	,
(	3236	)	,
(	3231	)	,
(	3226	)	,
(	3221	)	,
(	3216	)	,
(	3211	)	,
(	3207	)	,
(	3202	)	,
(	3197	)	,
(	3192	)	,
(	3187	)	,
(	3182	)	,
(	3178	)	,
(	3173	)	,
(	3168	)	,
(	3163	)	,
(	3159	)	,
(	3154	)	,
(	3149	)	,
(	3144	)	,
(	3139	)	,
(	3135	)	,
(	3130	)	,
(	3125	)	,
(	3121	)	,
(	3116	)	,
(	3111	)	,
(	3106	)	,
(	3102	)	,
(	3097	)	,
(	3092	)	,
(	3088	)	,
(	3083	)	,
(	3078	)	,
(	3074	)	,
(	3069	)	,
(	3064	)	,
(	3060	)	,
(	3055	)	,
(	3050	)	,
(	3046	)	,
(	3041	)	,
(	3036	)	,
(	3032	)	,
(	3027	)	,
(	3023	)	,
(	3018	)	,
(	3013	)	,
(	3009	)	,
(	3004	)	,
(	3000	)	,
(	2995	)	,
(	2990	)	,
(	2986	)	,
(	2981	)	,
(	2977	)	,
(	2972	)	,
(	2968	)	,
(	2963	)	,
(	2959	)	,
(	2954	)	,
(	2950	)	,
(	2945	)	,
(	2941	)	,
(	2936	)	,
(	2932	)	,
(	2927	)	,
(	2923	)	,
(	2918	)	,
(	2914	)	,
(	2909	)	,
(	2905	)	,
(	2900	)	,
(	2896	)	,
(	2892	)	,
(	2887	)	,
(	2883	)	,
(	2878	)	,
(	2874	)	,
(	2869	)	,
(	2865	)	,
(	2861	)	,
(	2856	)	,
(	2852	)	,
(	2848	)	,
(	2843	)	,
(	2839	)	,
(	2834	)	,
(	2830	)	,
(	2826	)	,
(	2821	)	,
(	2817	)	,
(	2813	)	,
(	2808	)	,
(	2804	)	,
(	2800	)	,
(	2795	)	,
(	2791	)	,
(	2787	)	,
(	2783	)	,
(	2778	)	,
(	2774	)	,
(	2770	)	,
(	2765	)	,
(	2761	)	,
(	2757	)	,
(	2753	)	,
(	2748	)	,
(	2744	)	,
(	2740	)	,
(	2736	)	,
(	2732	)	,
(	2727	)	,
(	2723	)	,
(	2719	)	,
(	2715	)	,
(	2711	)	,
(	2706	)	,
(	2702	)	,
(	2698	)	,
(	2694	)	,
(	2690	)	,
(	2685	)	,
(	2681	)	,
(	2677	)	,
(	2673	)	,
(	2669	)	,
(	2665	)	,
(	2661	)	,
(	2657	)	,
(	2652	)	,
(	2648	)	,
(	2644	)	,
(	2640	)	,
(	2636	)	,
(	2632	)	,
(	2628	)	,
(	2624	)	,
(	2620	)	,
(	2616	)	,
(	2612	)	,
(	2607	)	,
(	2603	)	,
(	2599	)	,
(	2595	)	,
(	2591	)	,
(	2587	)	,
(	2583	)	,
(	2579	)	,
(	2575	)	,
(	2571	)	,
(	2567	)	,
(	2563	)	,
(	2559	)	,
(	2555	)	,
(	2551	)	,
(	2547	)	,
(	2543	)	,
(	2539	)	,
(	2535	)	,
(	2532	)	,
(	2528	)	,
(	2524	)	,
(	2520	)	,
(	2516	)	,
(	2512	)	,
(	2508	)	,
(	2504	)	,
(	2500	)	,
(	2496	)	,
(	2492	)	,
(	2488	)	,
(	2485	)	,
(	2481	)	,
(	2477	)	,
(	2473	)	,
(	2469	)	,
(	2465	)	,
(	2461	)	,
(	2457	)	,
(	2454	)	,
(	2450	)	,
(	2446	)	,
(	2442	)	,
(	2438	)	,
(	2435	)	,
(	2431	)	,
(	2427	)	,
(	2423	)	,
(	2419	)	,
(	2416	)	,
(	2412	)	,
(	2408	)	,
(	2404	)	,
(	2400	)	,
(	2397	)	,
(	2393	)	,
(	2389	)	,
(	2385	)	,
(	2382	)	,
(	2378	)	,
(	2374	)	,
(	2370	)	,
(	2367	)	,
(	2363	)	,
(	2359	)	,
(	2356	)	,
(	2352	)	,
(	2348	)	,
(	2345	)	,
(	2341	)	,
(	2337	)	,
(	2334	)	,
(	2330	)	,
(	2326	)	,
(	2323	)	,
(	2319	)	,
(	2315	)	,
(	2312	)	,
(	2308	)	,
(	2304	)	,
(	2301	)	,
(	2297	)	,
(	2293	)	,
(	2290	)	,
(	2286	)	,
(	2283	)	,
(	2279	)	,
(	2275	)	,
(	2272	)	,
(	2268	)	,
(	2265	)	,
(	2261	)	,
(	2258	)	,
(	2254	)	,
(	2250	)	,
(	2247	)	,
(	2243	)	,
(	2240	)	,
(	2236	)	,
(	2233	)	,
(	2229	)	,
(	2226	)	,
(	2222	)	,
(	2219	)	,
(	2215	)	,
(	2212	)	,
(	2208	)	,
(	2205	)	,
(	2201	)	,
(	2198	)	,
(	2194	)	,
(	2191	)	,
(	2187	)	,
(	2184	)	,
(	2180	)	,
(	2177	)	,
(	2174	)	,
(	2170	)	,
(	2167	)	,
(	2163	)	,
(	2160	)	,
(	2156	)	,
(	2153	)	,
(	2150	)	,
(	2146	)	,
(	2143	)	,
(	2139	)	,
(	2136	)	,
(	2133	)	,
(	2129	)	,
(	2126	)	,
(	2123	)	,
(	2119	)	,
(	2116	)	,
(	2112	)	,
(	2109	)	,
(	2106	)	,
(	2102	)	,
(	2099	)	,
(	2096	)	,
(	2092	)	,
(	2089	)	,
(	2086	)	,
(	2083	)	,
(	2079	)	,
(	2076	)	,
(	2073	)	,
(	2069	)	,
(	2066	)	,
(	2063	)	,
(	2060	)	,
(	2056	)	,
(	2053	)	,
(	2050	)	,
(	2046	)	,
(	2043	)	,
(	2040	)	,
(	2037	)	,
(	2034	)	,
(	2030	)	,
(	2027	)	,
(	2024	)	,
(	2021	)	,
(	2017	)	,
(	2014	)	,
(	2011	)	,
(	2008	)	,
(	2005	)	,
(	2001	)	,
(	1998	)	,
(	1995	)	,
(	1992	)	,
(	1989	)	,
(	1986	)	,
(	1982	)	,
(	1979	)	,
(	1976	)	,
(	1973	)	,
(	1970	)	,
(	1967	)	,
(	1964	)	,
(	1960	)	,
(	1957	)	,
(	1954	)	,
(	1951	)	,
(	1948	)	,
(	1945	)	,
(	1942	)	,
(	1939	)	,
(	1936	)	,
(	1933	)	,
(	1929	)	,
(	1926	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1899	)	,
(	1896	)	,
(	1893	)	,
(	1890	)	,
(	1887	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1875	)	,
(	1872	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1857	)	,
(	1854	)	,
(	1851	)	,
(	1848	)	,
(	1845	)	,
(	1842	)	,
(	1839	)	,
(	1836	)	,
(	1833	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1765	)	,
(	1762	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1751	)	,
(	1748	)	,
(	1745	)	,
(	1742	)	,
(	1739	)	,
(	1737	)	,
(	1734	)	,
(	1731	)	,
(	1728	)	,
(	1726	)	,
(	1723	)	,
(	1720	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1709	)	,
(	1706	)	,
(	1704	)	,
(	1701	)	,
(	1698	)	,
(	1696	)	,
(	1693	)	,
(	1690	)	,
(	1687	)	,
(	1685	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1671	)	,
(	1669	)	,
(	1666	)	,
(	1663	)	,
(	1661	)	,
(	1658	)	,
(	1655	)	,
(	1653	)	,
(	1650	)	,
(	1648	)	,
(	1645	)	,
(	1642	)	,
(	1640	)	,
(	1637	)	,
(	1635	)	,
(	1632	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1619	)	,
(	1616	)	,
(	1614	)	,
(	1611	)	,
(	1609	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1598	)	,
(	1596	)	,
(	1593	)	,
(	1591	)	,
(	1588	)	,
(	1586	)	,
(	1583	)	,
(	1581	)	,
(	1578	)	,
(	1576	)	,
(	1573	)	,
(	1571	)	,
(	1568	)	,
(	1566	)	,
(	1563	)	,
(	1561	)	,
(	1558	)	,
(	1556	)	,
(	1553	)	,
(	1551	)	,
(	1548	)	,
(	1546	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1536	)	,
(	1534	)	,
(	1531	)	,
(	1529	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1519	)	,
(	1517	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1507	)	,
(	1505	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1495	)	,
(	1493	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1462	)	,
(	1460	)	,
(	1458	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1439	)	,
(	1437	)	,
(	1435	)	,
(	1433	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1382	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1349	)	,
(	1347	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1339	)	,
(	1337	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1328	)	,
(	1326	)	,
(	1324	)	,
(	1322	)	,
(	1320	)	,
(	1318	)	,
(	1316	)	,
(	1314	)	,
(	1312	)	,
(	1310	)	,
(	1308	)	,
(	1306	)	,
(	1304	)	,
(	1302	)	,
(	1300	)	,
(	1298	)	,
(	1296	)	,
(	1294	)	,
(	1292	)	,
(	1290	)	,
(	1288	)	,
(	1286	)	,
(	1284	)	,
(	1282	)	,
(	1280	)	,
(	1278	)	,
(	1276	)	,
(	1274	)	,
(	1272	)	,
(	1270	)	,
(	1268	)	,
(	1266	)	,
(	1264	)	,
(	1262	)	,
(	1260	)	,
(	1258	)	,
(	1256	)	,
(	1254	)	,
(	1252	)	,
(	1250	)	,
(	1248	)	,
(	1246	)	,
(	1244	)	,
(	1243	)	,
(	1241	)	,
(	1239	)	,
(	1237	)	,
(	1235	)	,
(	1233	)	,
(	1231	)	,
(	1229	)	,
(	1227	)	,
(	1225	)	,
(	1224	)	,
(	1222	)	,
(	1220	)	,
(	1218	)	,
(	1216	)	,
(	1214	)	,
(	1212	)	,
(	1210	)	,
(	1209	)	,
(	1207	)	,
(	1205	)	,
(	1203	)	,
(	1201	)	,
(	1199	)	,
(	1198	)	,
(	1196	)	,
(	1194	)	,
(	1192	)	,
(	1190	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1183	)	,
(	1181	)	,
(	1179	)	,
(	1178	)	,
(	1176	)	,
(	1174	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1160	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1151	)	,
(	1149	)	,
(	1148	)	,
(	1146	)	,
(	1144	)	,
(	1142	)	,
(	1141	)	,
(	1139	)	,
(	1137	)	,
(	1135	)	,
(	1134	)	,
(	1132	)	,
(	1130	)	,
(	1129	)	,
(	1127	)	,
(	1125	)	,
(	1124	)	,
(	1122	)	,
(	1120	)	,
(	1118	)	,
(	1117	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1110	)	,
(	1108	)	,
(	1107	)	,
(	1105	)	,
(	1104	)	,
(	1102	)	,
(	1100	)	,
(	1099	)	,
(	1097	)	,
(	1095	)	,
(	1094	)	,
(	1092	)	,
(	1090	)	,
(	1089	)	,
(	1087	)	,
(	1086	)	,
(	1084	)	,
(	1082	)	,
(	1081	)	,
(	1079	)	,
(	1078	)	,
(	1076	)	,
(	1074	)	,
(	1073	)	,
(	1071	)	,
(	1070	)	,
(	1068	)	,
(	1066	)	,
(	1065	)	,
(	1063	)	,
(	1062	)	,
(	1060	)	,
(	1059	)	,
(	1057	)	,
(	1055	)	,
(	1054	)	,
(	1052	)	,
(	1051	)	,
(	1049	)	,
(	1048	)	,
(	1046	)	,
(	1045	)	,
(	1043	)	,
(	1042	)	,
(	1040	)	,
(	1039	)	,
(	1037	)	,
(	1036	)	,
(	1034	)	,
(	1033	)	,
(	1031	)	,
(	1030	)	,
(	1028	)	,
(	1027	)	,
(	1025	)	,
(	1024	)	,
(	1022	)	,
(	1021	)	,
(	1019	)	,
(	1018	)	,
(	1016	)	,
(	1015	)	,
(	1013	)	,
(	1012	)	,
(	1010	)	,
(	1009	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1003	)	,
(	1002	)	,
(	1000	)	,
(	999	)	,
(	997	)	,
(	996	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	990	)	,
(	989	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	983	)	,
(	982	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	976	)	,
(	975	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	965	)	,
(	964	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	327	)	,
(	327	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	319	)	,
(	319	)	,
(	318	)	,
(	317	)	,
(	317	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	313	)	,
(	312	)	,
(	312	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	308	)	,
(	307	)	,
(	307	)	,
(	306	)	,
(	305	)	,
(	305	)	,
(	304	)	,
(	303	)	,
(	302	)	,
(	302	)	,
(	301	)	,
(	300	)	,
(	300	)	,
(	299	)	,
(	298	)	,
(	297	)	,
(	297	)	,
(	296	)	,
(	295	)	,
(	294	)	,
(	294	)	,
(	293	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	286	)	,
(	285	)	,
(	285	)	,
(	284	)	,
(	283	)	,
(	282	)	,
(	281	)	,
(	281	)	,
(	280	)	,
(	279	)	,
(	278	)	,
(	278	)	,
(	277	)	,
(	276	)	,
(	275	)	,
(	274	)	,
(	274	)	,
(	273	)	,
(	272	)	,
(	271	)	,
(	270	)	,
(	270	)	,
(	269	)	,
(	268	)	,
(	267	)	,
(	266	)	,
(	266	)	,
(	265	)	,
(	264	)	,
(	263	)	,
(	262	)	,
(	262	)	,
(	261	)	,
(	260	)	,
(	259	)	,
(	258	)	,
(	257	)	,
(	257	)	,
(	256	)	,
(	255	)	,
(	254	)	,
(	253	)	,
(	252	)	,
(	252	)	,
(	251	)	,
(	250	)	,
(	249	)	,
(	248	)	,
(	247	)	,
(	246	)	,
(	246	)	,
(	245	)	,
(	244	)	,
(	243	)	,
(	242	)	,
(	241	)	,
(	240	)	,
(	240	)	,
(	239	)	,
(	238	)	,
(	237	)	,
(	236	)	,
(	235	)	,
(	234	)	,
(	233	)	,
(	233	)	,
(	232	)	,
(	231	)	,
(	230	)	,
(	229	)	,
(	228	)	,
(	227	)	,
(	226	)	,
(	225	)	,
(	225	)	,
(	224	)	,
(	223	)	,
(	222	)	,
(	221	)	,
(	220	)	,
(	219	)	,
(	218	)	,
(	217	)	,
(	216	)	,
(	215	)	,
(	215	)	,
(	214	)	,
(	213	)	,
(	212	)	,
(	211	)	,
(	210	)	,
(	209	)	,
(	208	)	,
(	207	)	,
(	206	)	,
(	205	)	,
(	204	)	,
(	203	)	,
(	202	)	,
(	201	)	,
(	200	)	,
(	200	)	,
(	199	)	,
(	198	)	,
(	197	)	,
(	196	)	,
(	195	)	,
(	194	)	,
(	193	)	,
(	192	)	,
(	191	)	,
(	190	)	,
(	189	)	,
(	188	)	,
(	187	)	,
(	186	)	,
(	185	)	,
(	184	)	,
(	183	)	,
(	182	)	,
(	181	)	,
(	180	)	,
(	179	)	,
(	178	)	,
(	177	)	,
(	176	)	,
(	175	)	,
(	174	)	,
(	173	)	,
(	172	)	,
(	171	)	,
(	170	)	,
(	169	)	,
(	168	)	,
(	167	)	,
(	166	)	,
(	165	)	,
(	164	)	,
(	163	)	,
(	162	)	,
(	161	)	,
(	160	)	,
(	159	)	,
(	158	)	,
(	157	)	,
(	156	)	,
(	155	)	,
(	153	)	,
(	152	)	,
(	151	)	,
(	150	)	,
(	149	)	,
(	148	)	,
(	147	)	,
(	146	)	,
(	145	)	,
(	144	)	,
(	143	)	,
(	142	)	,
(	141	)	,
(	140	)	,
(	139	)	,
(	138	)	,
(	136	)	,
(	135	)	,
(	134	)	,
(	133	)	,
(	132	)	,
(	131	)	,
(	130	)	,
(	129	)	,
(	128	)	,
(	127	)	,
(	126	)	,
(	124	)	,
(	123	)	,
(	122	)	,
(	121	)	,
(	120	)	,
(	119	)	,
(	118	)	,
(	117	)	,
(	116	)	,
(	114	)	,
(	113	)	,
(	112	)	,
(	111	)	,
(	110	)	,
(	109	)	,
(	108	)	,
(	107	)	,
(	105	)	,
(	104	)	,
(	103	)	,
(	102	)	,
(	101	)	,
(	100	)	,
(	99	)	,
(	97	)	,
(	96	)	,
(	95	)	,
(	94	)	,
(	93	)	,
(	92	)	,
(	90	)	,
(	89	)	,
(	88	)	,
(	87	)	,
(	86	)	,
(	85	)	,
(	83	)	,
(	82	)	,
(	81	)	,
(	80	)	,
(	79	)	,
(	77	)	,
(	76	)	,
(	75	)	,
(	74	)	,
(	73	)	,
(	71	)	,
(	70	)	,
(	69	)	,
(	68	)	,
(	67	)	,
(	65	)	,
(	64	)	,
(	63	)	,
(	62	)	,
(	60	)	,
(	59	)	,
(	58	)	,
(	57	)	,
(	56	)	,
(	54	)	,
(	53	)	,
(	52	)	,
(	51	)	,
(	49	)	,
(	48	)	,
(	47	)	,
(	46	)	,
(	44	)	,
(	43	)	,
(	42	)	,
(	41	)	,
(	39	)	,
(	38	)	,
(	37	)	,
(	36	)	,
(	34	)	,
(	33	)	,
(	32	)	,
(	30	)	,
(	29	)	,
(	28	)	,
(	27	)	,
(	25	)	,
(	24	)	,
(	23	)	,
(	21	)	,
(	20	)	,
(	19	)	,
(	18	)	,
(	16	)	,
(	15	)	,
(	14	)	,
(	12	)	,
(	11	)	,
(	10	)	,
(	8	)	,
(	7	)	,
(	6	)	,
(	4	)	,
(	3	)	,
(	2	)	,
(	1	)	,
(	-1	)	,
(	-2	)	,
(	-3	)	,
(	-5	)	,
(	-6	)	,
(	-8	)	,
(	-9	)	,
(	-10	)	,
(	-12	)	,
(	-13	)	,
(	-14	)	,
(	-16	)	,
(	-17	)	,
(	-18	)	,
(	-20	)	,
(	-21	)	,
(	-22	)	,
(	-24	)	,
(	-25	)	,
(	-27	)	,
(	-28	)	,
(	-29	)	,
(	-31	)	,
(	-32	)	,
(	-33	)	,
(	-35	)	,
(	-36	)	,
(	-38	)	,
(	-39	)	,
(	-40	)	,
(	-42	)	,
(	-43	)	,
(	-45	)	,
(	-46	)	,
(	-47	)	,
(	-49	)	,
(	-50	)	,
(	-52	)	,
(	-53	)	,
(	-55	)	,
(	-56	)	,
(	-57	)	,
(	-59	)	,
(	-60	)	,
(	-62	)	,
(	-63	)	,
(	-65	)	,
(	-66	)	,
(	-67	)	,
(	-69	)	,
(	-70	)	,
(	-72	)	,
(	-73	)	,
(	-75	)	,
(	-76	)	,
(	-78	)	,
(	-79	)	,
(	-81	)	,
(	-82	)	,
(	-83	)	,
(	-85	)	,
(	-86	)	,
(	-88	)	,
(	-89	)	,
(	-91	)	,
(	-92	)	,
(	-94	)	,
(	-95	)	,
(	-97	)	,
(	-98	)	,
(	-100	)	,
(	-101	)	,
(	-103	)	,
(	-104	)	,
(	-106	)	,
(	-107	)	,
(	-109	)	,
(	-110	)	,
(	-112	)	,
(	-113	)	,
(	-115	)	,
(	-116	)	,
(	-118	)	,
(	-120	)	,
(	-121	)	,
(	-123	)	,
(	-124	)	,
(	-126	)	,
(	-127	)	,
(	-129	)	,
(	-130	)	,
(	-132	)	,
(	-133	)	,
(	-135	)	,
(	-136	)	,
(	-138	)	,
(	-140	)	,
(	-141	)	,
(	-143	)	,
(	-144	)	,
(	-146	)	,
(	-147	)	,
(	-149	)	,
(	-151	)	,
(	-152	)	,
(	-154	)	,
(	-155	)	,
(	-157	)	,
(	-159	)	,
(	-160	)	,
(	-162	)	,
(	-163	)	,
(	-165	)	,
(	-167	)	,
(	-168	)	,
(	-170	)	,
(	-171	)	,
(	-173	)	,
(	-175	)	,
(	-176	)	,
(	-178	)	,
(	-179	)	,
(	-181	)	,
(	-183	)	,
(	-184	)	,
(	-186	)	,
(	-188	)	,
(	-189	)	,
(	-191	)	,
(	-193	)	,
(	-194	)	,
(	-196	)	,
(	-197	)	,
(	-199	)	,
(	-201	)	,
(	-202	)	,
(	-204	)	,
(	-206	)	,
(	-207	)	,
(	-209	)	,
(	-211	)	,
(	-212	)	,
(	-214	)	,
(	-216	)	,
(	-217	)	,
(	-219	)	,
(	-221	)	,
(	-223	)	,
(	-224	)	,
(	-226	)	,
(	-228	)	,
(	-229	)	,
(	-231	)	,
(	-233	)	,
(	-234	)	,
(	-236	)	,
(	-238	)	,
(	-240	)	,
(	-241	)	,
(	-243	)	,
(	-245	)	,
(	-246	)	,
(	-248	)	,
(	-250	)	,
(	-252	)	,
(	-253	)	,
(	-255	)	,
(	-257	)	,
(	-259	)	,
(	-260	)	,
(	-262	)	,
(	-264	)	,
(	-266	)	,
(	-267	)	,
(	-269	)	,
(	-271	)	,
(	-273	)	,
(	-274	)	,
(	-276	)	,
(	-278	)	,
(	-280	)	,
(	-282	)	,
(	-283	)	,
(	-285	)	,
(	-287	)	,
(	-289	)	,
(	-290	)	,
(	-292	)	,
(	-294	)	,
(	-296	)	,
(	-298	)	,
(	-299	)	,
(	-301	)	,
(	-303	)	,
(	-305	)	,
(	-307	)	,
(	-309	)	,
(	-310	)	,
(	-312	)	,
(	-314	)	,
(	-316	)	,
(	-318	)	,
(	-319	)	,
(	-321	)	,
(	-323	)	,
(	-325	)	,
(	-327	)	,
(	-329	)	,
(	-331	)	,
(	-332	)	,
(	-334	)	,
(	-336	)	,
(	-338	)	,
(	-340	)	,
(	-342	)	,
(	-344	)	,
(	-345	)	,
(	-347	)	,
(	-349	)	,
(	-351	)	,
(	-353	)	,
(	-355	)	,
(	-357	)	,
(	-359	)	,
(	-360	)	,
(	-362	)	,
(	-364	)	,
(	-366	)	,
(	-368	)	,
(	-370	)	,
(	-372	)	,
(	-374	)	,
(	-376	)	,
(	-378	)	,
(	-380	)	,
(	-381	)	,
(	-383	)	,
(	-385	)	,
(	-387	)	,
(	-389	)	,
(	-391	)	,
(	-393	)	,
(	-395	)	,
(	-397	)	,
(	-399	)	,
(	-401	)	,
(	-403	)	,
(	-405	)	,
(	-407	)	,
(	-409	)	,
(	-411	)	,
(	-413	)	,
(	-415	)	,
(	-416	)	,
(	-418	)	,
(	-420	)	,
(	-422	)	,
(	-424	)	,
(	-426	)	,
(	-428	)	,
(	-430	)	,
(	-432	)	,
(	-434	)	,
(	-436	)	,
(	-438	)	,
(	-440	)	,
(	-442	)	,
(	-444	)	,
(	-446	)	,
(	-448	)	,
(	-450	)	,
(	-452	)	,
(	-454	)	,
(	-456	)	,
(	-458	)	,
(	-461	)	,
(	-463	)	,
(	-465	)	,
(	-467	)	,
(	-469	)	,
(	-471	)	,
(	-473	)	,
(	-475	)	,
(	-477	)	,
(	-479	)	,
(	-481	)	,
(	-483	)	,
(	-485	)	,
(	-487	)	,
(	-489	)	,
(	-491	)	,
(	-493	)	,
(	-495	)	,
(	-498	)	,
(	-500	)	,
(	-502	)	,
(	-504	)	,
(	-506	)	,
(	-508	)	,
(	-510	)	,
(	-512	)	,
(	-514	)	,
(	-516	)	,
(	-518	)	,
(	-521	)	,
(	-523	)	,
(	-525	)	,
(	-527	)	,
(	-529	)	,
(	-531	)	,
(	-533	)	,
(	-535	)	,
(	-538	)	,
(	-540	)	,
(	-542	)	,
(	-544	)	,
(	-546	)	,
(	-548	)	,
(	-550	)	,
(	-553	)	,
(	-555	)	,
(	-557	)	,
(	-559	)	,
(	-561	)	,
(	-563	)	,
(	-566	)	,
(	-568	)	,
(	-570	)	,
(	-572	)	,
(	-574	)	,
(	-576	)	,
(	-579	)	,
(	-581	)	,
(	-583	)	,
(	-585	)	,
(	-587	)	,
(	-590	)	,
(	-592	)	,
(	-594	)	,
(	-596	)	,
(	-598	)	,
(	-601	)	,
(	-603	)	,
(	-605	)	,
(	-607	)	,
(	-610	)	,
(	-612	)	,
(	-614	)	,
(	-616	)	,
(	-619	)	,
(	-621	)	,
(	-623	)	,
(	-625	)	,
(	-628	)	,
(	-630	)	,
(	-632	)	,
(	-634	)	,
(	-637	)	,
(	-639	)	,
(	-641	)	,
(	-643	)	,
(	-646	)	,
(	-648	)	,
(	-650	)	,
(	-652	)	,
(	-655	)	,
(	-657	)	,
(	-659	)	,
(	-662	)	,
(	-664	)	,
(	-666	)	,
(	-669	)	,
(	-671	)	,
(	-673	)	,
(	-675	)	,
(	-678	)	,
(	-680	)	,
(	-682	)	,
(	-685	)	,
(	-687	)	,
(	-689	)	,
(	-692	)	,
(	-694	)	,
(	-696	)	,
(	-699	)	,
(	-701	)	,
(	-703	)	,
(	-706	)	,
(	-708	)	,
(	-710	)	,
(	-713	)	,
(	-715	)	,
(	-718	)	,
(	-720	)	,
(	-722	)	,
(	-725	)	,
(	-727	)	,
(	-729	)	,
(	-732	)	,
(	-734	)	,
(	-737	)	,
(	-739	)	,
(	-741	)	,
(	-744	)	,
(	-746	)	,
(	-749	)	,
(	-751	)	,
(	-753	)	,
(	-756	)	,
(	-758	)	,
(	-761	)	,
(	-763	)	,
(	-765	)	,
(	-768	)	,
(	-770	)	,
(	-773	)	,
(	-775	)	,
(	-778	)	,
(	-780	)	,
(	-782	)	,
(	-785	)	,
(	-787	)	,
(	-790	)	,
(	-792	)	,
(	-795	)	,
(	-797	)	,
(	-800	)	,
(	-802	)	,
(	-805	)	,
(	-807	)	,
(	-810	)	,
(	-812	)	,
(	-815	)	,
(	-817	)	,
(	-819	)	,
(	-822	)	,
(	-824	)	,
(	-827	)	,
(	-829	)	,
(	-832	)	,
(	-834	)	,
(	-837	)	,
(	-839	)	,
(	-842	)	,
(	-845	)	,
(	-847	)	,
(	-850	)	,
(	-852	)	,
(	-855	)	,
(	-857	)	,
(	-860	)	,
(	-862	)	,
(	-865	)	,
(	-867	)	,
(	-870	)	,
(	-872	)	,
(	-875	)	,
(	-878	)	,
(	-880	)	,
(	-883	)	,
(	-885	)	,
(	-888	)	,
(	-890	)	,
(	-893	)	,
(	-896	)	,
(	-898	)	,
(	-901	)	,
(	-903	)	,
(	-906	)	,
(	-908	)	,
(	-911	)	,
(	-914	)	,
(	-916	)	,
(	-919	)	,
(	-921	)	,
(	-924	)	,
(	-927	)	,
(	-929	)	,
(	-932	)	,
(	-935	)	,
(	-937	)	,
(	-940	)	,
(	-942	)	,
(	-945	)	,
(	-948	)	,
(	-950	)	,
(	-953	)	,
(	-956	)	,
(	-958	)	,
(	-961	)	,
(	-964	)	,
(	-966	)	,
(	-969	)	,
(	-972	)	,
(	-974	)	,
(	-977	)	,
(	-980	)	,
(	-982	)	,
(	-985	)	,
(	-988	)	,
(	-990	)	,
(	-993	)	,
(	-996	)	,
(	-998	)	,
(	-1001	)	,
(	-1004	)	,
(	-1007	)	,
(	-1009	)	,
(	-1012	)	,
(	-1015	)	,
(	-1017	)	,
(	-1020	)	,
(	-1023	)	,
(	-1026	)	,
(	-1028	)	,
(	-1031	)	,
(	-1034	)	,
(	-1037	)	,
(	-1039	)	,
(	-1042	)	,
(	-1045	)	,
(	-1048	)	,
(	-1050	)	,
(	-1053	)	,
(	-1056	)	,
(	-1059	)	,
(	-1061	)	,
(	-1064	)	,
(	-1067	)	,
(	-1070	)	,
(	-1072	)	,
(	-1075	)	,
(	-1078	)	,
(	-1081	)	,
(	-1084	)	,
(	-1086	)	,
(	-1089	)	,
(	-1092	)	,
(	-1095	)	,
(	-1098	)	,
(	-1100	)	,
(	-1103	)	,
(	-1106	)	,
(	-1109	)	,
(	-1112	)	,
(	-1115	)	,
(	-1117	)	,
(	-1120	)	,
(	-1123	)	,
(	-1126	)	,
(	-1129	)	,
(	-1132	)	,
(	-1134	)	,
(	-1137	)	,
(	-1140	)	,
(	-1143	)	,
(	-1146	)	,
(	-1149	)	,
(	-1152	)	,
(	-1154	)	,
(	-1157	)	,
(	-1160	)	,
(	-1163	)	,
(	-1166	)	,
(	-1169	)	,
(	-1172	)	,
(	-1175	)	,
(	-1178	)	,
(	-1180	)	,
(	-1183	)	,
(	-1186	)	,
(	-1189	)	,
(	-1192	)	,
(	-1195	)	,
(	-1198	)	,
(	-1201	)	,
(	-1204	)	,
(	-1207	)	,
(	-1210	)	,
(	-1213	)	,
(	-1216	)	,
(	-1218	)	,
(	-1221	)	,
(	-1224	)	,
(	-1227	)	,
(	-1230	)	,
(	-1233	)	,
(	-1236	)	,
(	-1239	)	,
(	-1242	)	,
(	-1245	)	,
(	-1248	)	,
(	-1251	)	,
(	-1254	)	,
(	-1257	)	,
(	-1260	)	,
(	-1263	)	,
(	-1266	)	,
(	-1269	)	,
(	-1272	)	,
(	-1275	)	,
(	-1278	)	,
(	-1281	)	,
(	-1284	)	,
(	-1287	)	,
(	-1290	)	,
(	-1293	)	,
(	-1296	)	,
(	-1299	)	,
(	-1302	)	,
(	-1305	)	,
(	-1308	)	,
(	-1311	)	,
(	-1314	)	,
(	-1317	)	,
(	-1320	)	,
(	-1323	)	,
(	-1326	)	,
(	-1330	)	,
(	-1333	)	,
(	-1336	)	,
(	-1339	)	,
(	-1342	)	,
(	-1345	)	,
(	-1348	)	,
(	-1351	)	,
(	-1354	)	,
(	-1357	)	,
(	-1360	)	,
(	-1363	)	,
(	-1366	)	,
(	-1370	)	,
(	-1373	)	,
(	-1376	)	,
(	-1379	)	,
(	-1382	)	,
(	-1385	)	,
(	-1388	)	,
(	-1391	)	,
(	-1395	)	,
(	-1398	)	,
(	-1401	)	,
(	-1404	)	,
(	-1407	)	,
(	-1410	)	,
(	-1413	)	,
(	-1417	)	,
(	-1420	)	,
(	-1423	)	,
(	-1426	)	,
(	-1429	)	,
(	-1432	)	,
(	-1435	)	,
(	-1439	)	,
(	-1442	)	,
(	-1445	)	,
(	-1448	)	,
(	-1451	)	,
(	-1455	)	,
(	-1458	)	,
(	-1461	)	,
(	-1464	)	,
(	-1467	)	,
(	-1471	)	,
(	-1474	)	,
(	-1477	)	,
(	-1480	)	,
(	-1483	)	,
(	-1487	)	,
(	-1490	)	,
(	-1493	)	,
(	-1496	)	,
(	-1500	)	,
(	-1503	)	,
(	-1506	)	,
(	-1509	)	,
(	-1513	)	,
(	-1516	)	,
(	-1519	)	,
(	-1522	)	,
(	-1526	)	,
(	-1529	)	,
(	-1532	)	,
(	-1535	)	,
(	-1539	)	,
(	-1542	)	,
(	-1545	)	,
(	-1548	)	,
(	-1552	)	,
(	-1555	)	,
(	-1558	)	,
(	-1562	)	,
(	-1565	)	,
(	-1568	)	,
(	-1572	)	,
(	-1575	)	,
(	-1578	)	,
(	-1582	)	,
(	-1585	)	,
(	-1588	)	,
(	-1591	)	,
(	-1595	)	,
(	-1598	)	,
(	-1602	)	,
(	-1605	)	,
(	-1608	)	,
(	-1612	)	,
(	-1615	)	,
(	-1618	)	,
(	-1622	)	,
(	-1625	)	,
(	-1628	)	,
(	-1632	)	,
(	-1635	)	,
(	-1638	)	,
(	-1642	)	,
(	-1645	)	,
(	-1649	)	,
(	-1652	)	,
(	-1655	)	,
(	-1659	)	,
(	-1662	)	,
(	-1666	)	,
(	-1669	)	,
(	-1672	)	,
(	-1676	)	,
(	-1679	)	,
(	-1683	)	,
(	-1686	)	,
(	-1689	)	,
(	-1693	)	,
(	-1696	)	,
(	-1700	)	,
(	-1703	)	,
(	-1707	)	,
(	-1710	)	,
(	-1714	)	,
(	-1717	)	,
(	-1720	)	,
(	-1724	)	,
(	-1727	)	,
(	-1731	)	,
(	-1734	)	,
(	-1738	)	,
(	-1741	)	,
(	-1745	)	,
(	-1748	)	,
(	-1752	)	,
(	-1755	)	,
(	-1759	)	,
(	-1762	)	,
(	-1766	)	,
(	-1769	)	,
(	-1773	)	,
(	-1776	)	,
(	-1780	)	,
(	-1783	)	,
(	-1787	)	,
(	-1790	)	,
(	-1794	)	,
(	-1797	)	,
(	-1801	)	,
(	-1804	)	,
(	-1808	)	,
(	-1811	)	,
(	-1815	)	,
(	-1819	)	,
(	-1822	)	,
(	-1826	)	,
(	-1829	)	,
(	-1833	)	,
(	-1836	)	,
(	-1840	)	,
(	-1843	)	,
(	-1847	)	,
(	-1851	)	,
(	-1854	)	,
(	-1858	)	,
(	-1861	)	,
(	-1865	)	,
(	-1869	)	,
(	-1872	)	,
(	-1876	)	,
(	-1879	)	,
(	-1883	)	,
(	-1887	)	,
(	-1890	)	,
(	-1894	)	,
(	-1897	)	,
(	-1901	)	,
(	-1905	)	,
(	-1908	)	,
(	-1912	)	,
(	-1916	)	,
(	-1919	)	,
(	-1923	)	,
(	-1927	)	,
(	-1930	)	,
(	-1934	)	,
(	-1938	)	,
(	-1941	)	,
(	-1945	)	,
(	-1949	)	,
(	-1952	)	,
(	-1956	)	,
(	-1960	)	,
(	-1963	)	,
(	-1967	)	,
(	-1971	)	,
(	-1974	)	,
(	-1978	)	,
(	-1982	)	,
(	-1985	)	,
(	-1989	)	,
(	-1993	)	,
(	-1997	)	,
(	-2000	)	,
(	-2004	)	,
(	-2008	)	,
(	-2011	)	,
(	-2015	)	,
(	-2019	)	,
(	-2023	)	,
(	-2026	)	,
(	-2030	)	,
(	-2034	)	,
(	-2038	)	,
(	-2041	)	,
(	-2045	)	,
(	-2049	)	,
(	-2053	)	,
(	-2056	)	,
(	-2060	)	,
(	-2064	)	,
(	-2068	)	,
(	-2072	)	,
(	-2075	)	,
(	-2079	)	,
(	-2083	)	,
(	-2087	)	,
(	-2091	)	,
(	-2094	)	,
(	-2098	)	,
(	-2102	)	,
(	-2106	)	,
(	-2110	)	,
(	-2113	)	,
(	-2117	)	,
(	-2121	)	,
(	-2125	)	,
(	-2129	)	,
(	-2133	)	,
(	-2136	)	,
(	-2140	)	,
(	-2144	)	,
(	-2148	)	,
(	-2152	)	,
(	-2156	)	,
(	-2160	)	,
(	-2163	)	,
(	-2167	)	,
(	-2171	)	,
(	-2175	)	,
(	-2179	)	,
(	-2183	)	,
(	-2187	)	,
(	-2191	)	,
(	-2195	)	,
(	-2198	)	,
(	-2202	)	,
(	-2206	)	,
(	-2210	)	,
(	-2214	)	,
(	-2218	)	,
(	-2222	)	,
(	-2226	)	,
(	-2230	)	,
(	-2234	)	,
(	-2238	)	,
(	-2242	)	,
(	-2245	)	,
(	-2249	)	,
(	-2253	)	,
(	-2257	)	,
(	-2261	)	,
(	-2265	)	,
(	-2269	)	,
(	-2273	)	,
(	-2277	)	,
(	-2281	)	,
(	-2285	)	,
(	-2289	)	,
(	-2293	)	,
(	-2297	)	,
(	-2301	)	,
(	-2305	)	,
(	-2309	)	,
(	-2313	)	,
(	-2317	)	,
(	-2321	)	,
(	-2325	)	,
(	-2329	)	,
(	-2333	)	,
(	-2337	)	,
(	-2341	)	,
(	-2345	)	,
(	-2349	)	,
(	-2353	)	,
(	-2357	)	,
(	-2361	)	,
(	-2365	)	,
(	-2369	)	,
(	-2373	)	,
(	-2377	)	,
(	-2382	)	,
(	-2386	)	,
(	-2390	)	,
(	-2394	)	,
(	-2398	)	,
(	-2402	)	,
(	-2406	)	,
(	-2410	)	,
(	-2414	)	,
(	-2418	)	,
(	-2422	)	,
(	-2426	)	,
(	-2431	)	,
(	-2435	)	,
(	-2439	)	,
(	-2443	)	,
(	-2447	)	,
(	-2451	)	,
(	-2455	)	,
(	-2459	)	,
(	-2463	)	,
(	-2468	)	,
(	-2472	)	,
(	-2476	)	,
(	-2480	)	,
(	-2484	)	,
(	-2488	)	,
(	-2492	)	,
(	-2497	)	,
(	-2501	)	,
(	-2505	)	,
(	-2509	)	,
(	-2513	)	,
(	-2517	)	,
(	-2522	)	,
(	-2526	)	,
(	-2530	)	,
(	-2534	)	,
(	-2538	)	,
(	-2543	)	,
(	-2547	)	,
(	-2551	)	,
(	-2555	)	,
(	-2559	)	,
(	-2564	)	,
(	-2568	)	,
(	-2572	)	,
(	-2576	)	,
(	-2581	)	,
(	-2585	)	,
(	-2589	)	,
(	-2593	)	,
(	-2598	)	,
(	-2602	)	,
(	-2606	)	,
(	-2610	)	,
(	-2615	)	,
(	-2619	)	,
(	-2623	)	,
(	-2627	)	,
(	-2632	)	,
(	-2636	)	,
(	-2640	)	,
(	-2644	)	,
(	-2649	)	,
(	-2653	)	,
(	-2657	)	,
(	-2662	)	,
(	-2666	)	,
(	-2670	)	,
(	-2675	)	,
(	-2679	)	,
(	-2683	)	,
(	-2687	)	,
(	-2692	)	,
(	-2696	)	,
(	-2700	)	,
(	-2705	)	,
(	-2709	)	,
(	-2713	)	,
(	-2718	)	,
(	-2722	)	,
(	-2726	)	,
(	-2731	)	,
(	-2735	)	,
(	-2740	)	,
(	-2744	)	,
(	-2748	)	,
(	-2753	)	,
(	-2757	)	,
(	-2761	)	,
(	-2766	)	,
(	-2770	)	,
(	-2775	)	,
(	-2779	)	,
(	-2783	)	,
(	-2788	)	,
(	-2792	)	,
(	-2797	)	,
(	-2801	)	,
(	-2805	)	,
(	-2810	)	,
(	-2814	)	,
(	-2819	)	,
(	-2823	)	,
(	-2828	)	,
(	-2832	)	,
(	-2836	)	,
(	-2841	)	,
(	-2845	)	,
(	-2850	)	,
(	-2854	)	,
(	-2859	)	,
(	-2863	)	,
(	-2868	)	,
(	-2872	)	,
(	-2877	)	,
(	-2881	)	,
(	-2886	)	,
(	-2890	)	,
(	-2894	)	,
(	-2899	)	,
(	-2903	)	,
(	-2908	)	,
(	-2912	)	,
(	-2917	)	,
(	-2921	)	,
(	-2926	)	,
(	-2931	)	,
(	-2935	)	,
(	-2940	)	,
(	-2944	)	,
(	-2949	)	,
(	-2953	)	,
(	-2958	)	,
(	-2962	)	,
(	-2967	)	,
(	-2971	)	,
(	-2976	)	,
(	-2980	)	,
(	-2985	)	,
(	-2990	)	,
(	-2994	)	,
(	-2999	)	,
(	-3003	)	,
(	-3008	)	,
(	-3012	)	,
(	-3017	)	,
(	-3022	)	,
(	-3026	)	,
(	-3031	)	,
(	-3035	)	,
(	-3040	)	,
(	-3045	)	,
(	-3049	)	,
(	-3054	)	,
(	-3058	)	,
(	-3063	)	,
(	-3068	)	,
(	-3072	)	,
(	-3077	)	,
(	-3082	)	,
(	-3086	)	,
(	-3091	)	,
(	-3096	)	,
(	-3100	)	,
(	-3105	)	,
(	-3110	)	,
(	-3114	)	,
(	-3119	)	,
(	-3124	)	,
(	-3128	)	,
(	-3133	)	,
(	-3138	)	,
(	-3142	)	,
(	-3147	)	,
(	-3152	)	,
(	-3156	)	,
(	-3161	)	,
(	-3166	)	,
(	-3170	)	,
(	-3175	)	,
(	-3180	)	,
(	-3185	)	,
(	-3189	)	,
(	-3194	)	,
(	-3199	)	,
(	-3203	)	,
(	-3208	)	,
(	-3213	)	,
(	-3218	)	,
(	-3222	)	,
(	-3227	)	,
(	-3232	)	,
(	-3237	)	
);



end package LUT_pkg;
