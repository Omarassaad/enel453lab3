library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	7855	)	,
(	7837	)	,
(	7818	)	,
(	7800	)	,
(	7782	)	,
(	7764	)	,
(	7746	)	,
(	7728	)	,
(	7710	)	,
(	7692	)	,
(	7674	)	,
(	7656	)	,
(	7638	)	,
(	7620	)	,
(	7603	)	,
(	7585	)	,
(	7567	)	,
(	7550	)	,
(	7532	)	,
(	7514	)	,
(	7497	)	,
(	7479	)	,
(	7462	)	,
(	7444	)	,
(	7427	)	,
(	7410	)	,
(	7392	)	,
(	7375	)	,
(	7358	)	,
(	7341	)	,
(	7323	)	,
(	7306	)	,
(	7289	)	,
(	7272	)	,
(	7255	)	,
(	7238	)	,
(	7221	)	,
(	7204	)	,
(	7187	)	,
(	7171	)	,
(	7154	)	,
(	7137	)	,
(	7120	)	,
(	7104	)	,
(	7087	)	,
(	7070	)	,
(	7054	)	,
(	7037	)	,
(	7021	)	,
(	7004	)	,
(	6988	)	,
(	6971	)	,
(	6955	)	,
(	6939	)	,
(	6923	)	,
(	6906	)	,
(	6890	)	,
(	6874	)	,
(	6858	)	,
(	6842	)	,
(	6826	)	,
(	6810	)	,
(	6794	)	,
(	6778	)	,
(	6762	)	,
(	6746	)	,
(	6730	)	,
(	6714	)	,
(	6698	)	,
(	6683	)	,
(	6667	)	,
(	6651	)	,
(	6635	)	,
(	6620	)	,
(	6604	)	,
(	6589	)	,
(	6573	)	,
(	6558	)	,
(	6542	)	,
(	6527	)	,
(	6512	)	,
(	6496	)	,
(	6481	)	,
(	6466	)	,
(	6450	)	,
(	6435	)	,
(	6420	)	,
(	6405	)	,
(	6390	)	,
(	6375	)	,
(	6360	)	,
(	6345	)	,
(	6330	)	,
(	6315	)	,
(	6300	)	,
(	6285	)	,
(	6270	)	,
(	6256	)	,
(	6241	)	,
(	6226	)	,
(	6211	)	,
(	6197	)	,
(	6182	)	,
(	6167	)	,
(	6153	)	,
(	6138	)	,
(	6124	)	,
(	6109	)	,
(	6095	)	,
(	6081	)	,
(	6066	)	,
(	6052	)	,
(	6038	)	,
(	6023	)	,
(	6009	)	,
(	5995	)	,
(	5981	)	,
(	5967	)	,
(	5953	)	,
(	5939	)	,
(	5925	)	,
(	5911	)	,
(	5897	)	,
(	5883	)	,
(	5869	)	,
(	5855	)	,
(	5841	)	,
(	5827	)	,
(	5813	)	,
(	5800	)	,
(	5786	)	,
(	5772	)	,
(	5759	)	,
(	5745	)	,
(	5732	)	,
(	5718	)	,
(	5704	)	,
(	5691	)	,
(	5678	)	,
(	5664	)	,
(	5651	)	,
(	5637	)	,
(	5624	)	,
(	5611	)	,
(	5597	)	,
(	5584	)	,
(	5571	)	,
(	5558	)	,
(	5545	)	,
(	5532	)	,
(	5519	)	,
(	5505	)	,
(	5492	)	,
(	5479	)	,
(	5467	)	,
(	5454	)	,
(	5441	)	,
(	5428	)	,
(	5415	)	,
(	5402	)	,
(	5389	)	,
(	5377	)	,
(	5364	)	,
(	5351	)	,
(	5339	)	,
(	5326	)	,
(	5313	)	,
(	5301	)	,
(	5288	)	,
(	5276	)	,
(	5263	)	,
(	5251	)	,
(	5239	)	,
(	5226	)	,
(	5214	)	,
(	5201	)	,
(	5189	)	,
(	5177	)	,
(	5165	)	,
(	5152	)	,
(	5140	)	,
(	5128	)	,
(	5116	)	,
(	5104	)	,
(	5092	)	,
(	5080	)	,
(	5068	)	,
(	5056	)	,
(	5044	)	,
(	5032	)	,
(	5020	)	,
(	5008	)	,
(	4996	)	,
(	4985	)	,
(	4973	)	,
(	4961	)	,
(	4949	)	,
(	4938	)	,
(	4926	)	,
(	4914	)	,
(	4903	)	,
(	4891	)	,
(	4880	)	,
(	4868	)	,
(	4857	)	,
(	4845	)	,
(	4834	)	,
(	4822	)	,
(	4811	)	,
(	4800	)	,
(	4788	)	,
(	4777	)	,
(	4766	)	,
(	4755	)	,
(	4743	)	,
(	4732	)	,
(	4721	)	,
(	4710	)	,
(	4699	)	,
(	4688	)	,
(	4677	)	,
(	4666	)	,
(	4655	)	,
(	4644	)	,
(	4633	)	,
(	4622	)	,
(	4611	)	,
(	4600	)	,
(	4589	)	,
(	4579	)	,
(	4568	)	,
(	4557	)	,
(	4546	)	,
(	4536	)	,
(	4525	)	,
(	4514	)	,
(	4504	)	,
(	4493	)	,
(	4483	)	,
(	4472	)	,
(	4462	)	,
(	4451	)	,
(	4441	)	,
(	4430	)	,
(	4420	)	,
(	4410	)	,
(	4399	)	,
(	4389	)	,
(	4379	)	,
(	4368	)	,
(	4358	)	,
(	4348	)	,
(	4338	)	,
(	4328	)	,
(	4317	)	,
(	4307	)	,
(	4297	)	,
(	4287	)	,
(	4277	)	,
(	4267	)	,
(	4257	)	,
(	4247	)	,
(	4237	)	,
(	4227	)	,
(	4218	)	,
(	4208	)	,
(	4198	)	,
(	4188	)	,
(	4178	)	,
(	4169	)	,
(	4159	)	,
(	4149	)	,
(	4139	)	,
(	4130	)	,
(	4120	)	,
(	4111	)	,
(	4101	)	,
(	4091	)	,
(	4082	)	,
(	4072	)	,
(	4063	)	,
(	4053	)	,
(	4044	)	,
(	4035	)	,
(	4025	)	,
(	4016	)	,
(	4006	)	,
(	3997	)	,
(	3988	)	,
(	3979	)	,
(	3969	)	,
(	3960	)	,
(	3951	)	,
(	3942	)	,
(	3933	)	,
(	3924	)	,
(	3914	)	,
(	3905	)	,
(	3896	)	,
(	3887	)	,
(	3878	)	,
(	3869	)	,
(	3860	)	,
(	3851	)	,
(	3843	)	,
(	3834	)	,
(	3825	)	,
(	3816	)	,
(	3807	)	,
(	3798	)	,
(	3790	)	,
(	3781	)	,
(	3772	)	,
(	3764	)	,
(	3755	)	,
(	3746	)	,
(	3738	)	,
(	3729	)	,
(	3720	)	,
(	3712	)	,
(	3703	)	,
(	3695	)	,
(	3686	)	,
(	3678	)	,
(	3669	)	,
(	3661	)	,
(	3653	)	,
(	3644	)	,
(	3636	)	,
(	3628	)	,
(	3619	)	,
(	3611	)	,
(	3603	)	,
(	3594	)	,
(	3586	)	,
(	3578	)	,
(	3570	)	,
(	3562	)	,
(	3554	)	,
(	3545	)	,
(	3537	)	,
(	3529	)	,
(	3521	)	,
(	3513	)	,
(	3505	)	,
(	3497	)	,
(	3489	)	,
(	3481	)	,
(	3473	)	,
(	3466	)	,
(	3458	)	,
(	3450	)	,
(	3442	)	,
(	3434	)	,
(	3426	)	,
(	3419	)	,
(	3411	)	,
(	3403	)	,
(	3395	)	,
(	3388	)	,
(	3380	)	,
(	3373	)	,
(	3365	)	,
(	3357	)	,
(	3350	)	,
(	3342	)	,
(	3335	)	,
(	3327	)	,
(	3320	)	,
(	3312	)	,
(	3305	)	,
(	3297	)	,
(	3290	)	,
(	3283	)	,
(	3275	)	,
(	3268	)	,
(	3260	)	,
(	3253	)	,
(	3246	)	,
(	3239	)	,
(	3231	)	,
(	3224	)	,
(	3217	)	,
(	3210	)	,
(	3203	)	,
(	3195	)	,
(	3188	)	,
(	3181	)	,
(	3174	)	,
(	3167	)	,
(	3160	)	,
(	3153	)	,
(	3146	)	,
(	3139	)	,
(	3132	)	,
(	3125	)	,
(	3118	)	,
(	3111	)	,
(	3104	)	,
(	3098	)	,
(	3091	)	,
(	3084	)	,
(	3077	)	,
(	3070	)	,
(	3063	)	,
(	3057	)	,
(	3050	)	,
(	3043	)	,
(	3037	)	,
(	3030	)	,
(	3023	)	,
(	3017	)	,
(	3010	)	,
(	3003	)	,
(	2997	)	,
(	2990	)	,
(	2984	)	,
(	2977	)	,
(	2971	)	,
(	2964	)	,
(	2958	)	,
(	2951	)	,
(	2945	)	,
(	2938	)	,
(	2932	)	,
(	2926	)	,
(	2919	)	,
(	2913	)	,
(	2907	)	,
(	2900	)	,
(	2894	)	,
(	2888	)	,
(	2882	)	,
(	2875	)	,
(	2869	)	,
(	2863	)	,
(	2857	)	,
(	2851	)	,
(	2844	)	,
(	2838	)	,
(	2832	)	,
(	2826	)	,
(	2820	)	,
(	2814	)	,
(	2808	)	,
(	2802	)	,
(	2796	)	,
(	2790	)	,
(	2784	)	,
(	2778	)	,
(	2772	)	,
(	2766	)	,
(	2760	)	,
(	2754	)	,
(	2749	)	,
(	2743	)	,
(	2737	)	,
(	2731	)	,
(	2725	)	,
(	2720	)	,
(	2714	)	,
(	2708	)	,
(	2702	)	,
(	2697	)	,
(	2691	)	,
(	2685	)	,
(	2680	)	,
(	2674	)	,
(	2668	)	,
(	2663	)	,
(	2657	)	,
(	2652	)	,
(	2646	)	,
(	2640	)	,
(	2635	)	,
(	2629	)	,
(	2624	)	,
(	2618	)	,
(	2613	)	,
(	2608	)	,
(	2602	)	,
(	2597	)	,
(	2591	)	,
(	2586	)	,
(	2581	)	,
(	2575	)	,
(	2570	)	,
(	2565	)	,
(	2559	)	,
(	2554	)	,
(	2549	)	,
(	2544	)	,
(	2538	)	,
(	2533	)	,
(	2528	)	,
(	2523	)	,
(	2518	)	,
(	2512	)	,
(	2507	)	,
(	2502	)	,
(	2497	)	,
(	2492	)	,
(	2487	)	,
(	2482	)	,
(	2477	)	,
(	2472	)	,
(	2467	)	,
(	2462	)	,
(	2457	)	,
(	2452	)	,
(	2447	)	,
(	2442	)	,
(	2437	)	,
(	2432	)	,
(	2427	)	,
(	2422	)	,
(	2417	)	,
(	2413	)	,
(	2408	)	,
(	2403	)	,
(	2398	)	,
(	2393	)	,
(	2389	)	,
(	2384	)	,
(	2379	)	,
(	2374	)	,
(	2370	)	,
(	2365	)	,
(	2360	)	,
(	2355	)	,
(	2351	)	,
(	2346	)	,
(	2342	)	,
(	2337	)	,
(	2332	)	,
(	2328	)	,
(	2323	)	,
(	2319	)	,
(	2314	)	,
(	2310	)	,
(	2305	)	,
(	2301	)	,
(	2296	)	,
(	2292	)	,
(	2287	)	,
(	2283	)	,
(	2278	)	,
(	2274	)	,
(	2269	)	,
(	2265	)	,
(	2261	)	,
(	2256	)	,
(	2252	)	,
(	2248	)	,
(	2243	)	,
(	2239	)	,
(	2235	)	,
(	2230	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2201	)	,
(	2197	)	,
(	2192	)	,
(	2188	)	,
(	2184	)	,
(	2180	)	,
(	2176	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2100	)	,
(	2096	)	,
(	2093	)	,
(	2089	)	,
(	2085	)	,
(	2081	)	,
(	2077	)	,
(	2074	)	,
(	2070	)	,
(	2066	)	,
(	2062	)	,
(	2059	)	,
(	2055	)	,
(	2051	)	,
(	2047	)	,
(	2044	)	,
(	2040	)	,
(	2036	)	,
(	2033	)	,
(	2029	)	,
(	2026	)	,
(	2022	)	,
(	2018	)	,
(	2015	)	,
(	2011	)	,
(	2008	)	,
(	2004	)	,
(	2000	)	,
(	1997	)	,
(	1993	)	,
(	1990	)	,
(	1986	)	,
(	1983	)	,
(	1979	)	,
(	1976	)	,
(	1973	)	,
(	1969	)	,
(	1966	)	,
(	1962	)	,
(	1959	)	,
(	1955	)	,
(	1952	)	,
(	1949	)	,
(	1945	)	,
(	1942	)	,
(	1939	)	,
(	1935	)	,
(	1932	)	,
(	1929	)	,
(	1925	)	,
(	1922	)	,
(	1919	)	,
(	1916	)	,
(	1912	)	,
(	1909	)	,
(	1906	)	,
(	1903	)	,
(	1899	)	,
(	1896	)	,
(	1893	)	,
(	1890	)	,
(	1887	)	,
(	1883	)	,
(	1880	)	,
(	1877	)	,
(	1874	)	,
(	1871	)	,
(	1868	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1837	)	,
(	1834	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1763	)	,
(	1760	)	,
(	1757	)	,
(	1754	)	,
(	1752	)	,
(	1749	)	,
(	1746	)	,
(	1743	)	,
(	1741	)	,
(	1738	)	,
(	1735	)	,
(	1733	)	,
(	1730	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1720	)	,
(	1717	)	,
(	1714	)	,
(	1712	)	,
(	1709	)	,
(	1707	)	,
(	1704	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1694	)	,
(	1691	)	,
(	1689	)	,
(	1686	)	,
(	1684	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1672	)	,
(	1669	)	,
(	1667	)	,
(	1664	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1648	)	,
(	1645	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1631	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1620	)	,
(	1617	)	,
(	1615	)	,
(	1613	)	,
(	1611	)	,
(	1609	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1600	)	,
(	1597	)	,
(	1595	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1584	)	,
(	1582	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1572	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1563	)	,
(	1561	)	,
(	1559	)	,
(	1557	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1447	)	,
(	1445	)	,
(	1443	)	,
(	1441	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1430	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1417	)	,
(	1415	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1409	)	,
(	1407	)	,
(	1406	)	,
(	1404	)	,
(	1403	)	,
(	1401	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1389	)	,
(	1387	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1380	)	,
(	1378	)	,
(	1377	)	,
(	1375	)	,
(	1374	)	,
(	1372	)	,
(	1371	)	,
(	1370	)	,
(	1368	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1361	)	,
(	1359	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1347	)	,
(	1345	)	,
(	1344	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1324	)	,
(	1323	)	,
(	1321	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1307	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1302	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1297	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1292	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1282	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1275	)	,
(	1274	)	,
(	1273	)	,
(	1272	)	,
(	1270	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1266	)	,
(	1265	)	,
(	1263	)	,
(	1262	)	,
(	1261	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1249	)	,
(	1247	)	,
(	1246	)	,
(	1245	)	,
(	1244	)	,
(	1243	)	,
(	1242	)	,
(	1241	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	761	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	751	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	732	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	610	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	402	)	,
(	402	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	405	)	,
(	405	)	,
(	406	)	,
(	406	)	,
(	407	)	,
(	407	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	409	)	,
(	409	)	,
(	410	)	,
(	410	)	,
(	411	)	,
(	411	)	,
(	412	)	,
(	413	)	,
(	413	)	,
(	414	)	,
(	414	)	,
(	415	)	,
(	415	)	,
(	416	)	,
(	417	)	,
(	417	)	,
(	418	)	,
(	418	)	,
(	419	)	,
(	420	)	,
(	420	)	,
(	421	)	,
(	422	)	,
(	422	)	,
(	423	)	,
(	424	)	,
(	424	)	,
(	425	)	,
(	426	)	,
(	427	)	,
(	427	)	,
(	428	)	,
(	429	)	,
(	430	)	,
(	430	)	,
(	431	)	,
(	432	)	,
(	433	)	,
(	433	)	,
(	434	)	,
(	435	)	,
(	436	)	,
(	437	)	,
(	438	)	,
(	439	)	,
(	439	)	,
(	440	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	444	)	,
(	445	)	,
(	446	)	,
(	447	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	451	)	,
(	452	)	,
(	453	)	,
(	454	)	,
(	455	)	,
(	456	)	,
(	457	)	,
(	458	)	,
(	459	)	,
(	460	)	,
(	461	)	,
(	462	)	,
(	463	)	,
(	464	)	,
(	465	)	,
(	467	)	,
(	468	)	,
(	469	)	,
(	470	)	,
(	471	)	,
(	472	)	,
(	474	)	,
(	475	)	,
(	476	)	,
(	477	)	,
(	479	)	,
(	480	)	,
(	481	)	,
(	482	)	,
(	484	)	,
(	485	)	,
(	486	)	,
(	487	)	,
(	489	)	,
(	490	)	,
(	491	)	,
(	493	)	,
(	494	)	,
(	496	)	,
(	497	)	,
(	498	)	,
(	500	)	,
(	501	)	,
(	503	)	,
(	504	)	,
(	506	)	,
(	507	)	,
(	508	)	,
(	510	)	,
(	511	)	,
(	513	)	,
(	514	)	,
(	516	)	,
(	518	)	,
(	519	)	,
(	521	)	,
(	522	)	,
(	524	)	,
(	525	)	,
(	527	)	,
(	529	)	,
(	530	)	,
(	532	)	,
(	534	)	,
(	535	)	,
(	537	)	,
(	539	)	,
(	540	)	,
(	542	)	,
(	544	)	,
(	546	)	,
(	547	)	,
(	549	)	,
(	551	)	,
(	553	)	,
(	554	)	,
(	556	)	,
(	558	)	,
(	560	)	,
(	562	)	,
(	564	)	,
(	565	)	,
(	567	)	,
(	569	)	,
(	571	)	,
(	573	)	,
(	575	)	,
(	577	)	,
(	579	)	,
(	581	)	,
(	583	)	,
(	585	)	,
(	587	)	,
(	589	)	,
(	591	)	,
(	593	)	,
(	595	)	,
(	597	)	,
(	599	)	,
(	601	)	,
(	603	)	,
(	605	)	,
(	608	)	,
(	610	)	,
(	612	)	,
(	614	)	,
(	616	)	,
(	618	)	,
(	621	)	,
(	623	)	,
(	625	)	,
(	627	)	,
(	630	)	,
(	632	)	,
(	634	)	,
(	637	)	,
(	639	)	,
(	641	)	,
(	644	)	,
(	646	)	,
(	648	)	,
(	651	)	,
(	653	)	,
(	655	)	,
(	658	)	,
(	660	)	,
(	663	)	,
(	665	)	,
(	668	)	,
(	670	)	,
(	673	)	,
(	675	)	,
(	678	)	,
(	680	)	,
(	683	)	,
(	685	)	,
(	688	)	,
(	691	)	,
(	693	)	,
(	696	)	,
(	699	)	,
(	701	)	,
(	704	)	,
(	707	)	,
(	709	)	,
(	712	)	,
(	715	)	,
(	718	)	,
(	720	)	,
(	723	)	,
(	726	)	,
(	729	)	,
(	732	)	,
(	734	)	,
(	737	)	,
(	740	)	,
(	743	)	,
(	746	)	,
(	749	)	,
(	752	)	,
(	755	)	,
(	758	)	,
(	761	)	,
(	764	)	,
(	767	)	,
(	770	)	,
(	773	)	,
(	776	)	,
(	779	)	,
(	782	)	,
(	785	)	,
(	788	)	,
(	791	)	,
(	794	)	,
(	797	)	,
(	801	)	,
(	804	)	,
(	807	)	,
(	810	)	,
(	813	)	,
(	817	)	,
(	820	)	,
(	823	)	,
(	826	)	,
(	830	)	,
(	833	)	,
(	836	)	,
(	840	)	,
(	843	)	,
(	847	)	,
(	850	)	,
(	853	)	,
(	857	)	,
(	860	)	,
(	864	)	,
(	867	)	,
(	871	)	,
(	874	)	,
(	878	)	,
(	881	)	,
(	885	)	,
(	888	)	,
(	892	)	,
(	896	)	,
(	899	)	,
(	903	)	,
(	907	)	,
(	910	)	,
(	914	)	,
(	918	)	,
(	921	)	,
(	925	)	,
(	929	)	,
(	933	)	,
(	937	)	,
(	940	)	,
(	944	)	,
(	948	)	,
(	952	)	,
(	956	)	,
(	960	)	,
(	964	)	,
(	968	)	,
(	971	)	,
(	975	)	,
(	979	)	,
(	983	)	,
(	987	)	,
(	992	)	,
(	996	)	,
(	1000	)	,
(	1004	)	,
(	1008	)	,
(	1012	)	,
(	1016	)	,
(	1020	)	,
(	1024	)	,
(	1029	)	,
(	1033	)	,
(	1037	)	,
(	1041	)	,
(	1046	)	,
(	1050	)	,
(	1054	)	,
(	1059	)	,
(	1063	)	,
(	1067	)	,
(	1072	)	,
(	1076	)	,
(	1080	)	,
(	1085	)	,
(	1089	)	,
(	1094	)	,
(	1098	)	,
(	1103	)	,
(	1107	)	,
(	1112	)	,
(	1116	)	,
(	1121	)	,
(	1126	)	,
(	1130	)	,
(	1135	)	,
(	1140	)	,
(	1144	)	,
(	1149	)	,
(	1154	)	,
(	1158	)	,
(	1163	)	,
(	1168	)	,
(	1173	)	,
(	1177	)	,
(	1182	)	,
(	1187	)	,
(	1192	)	,
(	1197	)	,
(	1202	)	,
(	1207	)	,
(	1212	)	,
(	1217	)	,
(	1222	)	,
(	1227	)	,
(	1232	)	,
(	1237	)	,
(	1242	)	,
(	1247	)	,
(	1252	)	,
(	1257	)	,
(	1262	)	,
(	1267	)	,
(	1272	)	,
(	1278	)	,
(	1283	)	,
(	1288	)	,
(	1293	)	,
(	1299	)	,
(	1304	)	,
(	1309	)	,
(	1315	)	,
(	1320	)	,
(	1325	)	,
(	1331	)	,
(	1336	)	,
(	1342	)	,
(	1347	)	,
(	1353	)	,
(	1358	)	,
(	1364	)	,
(	1369	)	,
(	1375	)	,
(	1380	)	,
(	1386	)	,
(	1392	)	,
(	1397	)	,
(	1403	)	,
(	1409	)	,
(	1414	)	,
(	1420	)	,
(	1426	)	,
(	1431	)	,
(	1437	)	,
(	1443	)	,
(	1449	)	,
(	1455	)	,
(	1461	)	,
(	1467	)	,
(	1472	)	,
(	1478	)	,
(	1484	)	,
(	1490	)	,
(	1496	)	,
(	1502	)	,
(	1508	)	,
(	1515	)	,
(	1521	)	,
(	1527	)	,
(	1533	)	,
(	1539	)	,
(	1545	)	,
(	1551	)	,
(	1558	)	,
(	1564	)	,
(	1570	)	,
(	1576	)	,
(	1583	)	,
(	1589	)	,
(	1595	)	,
(	1602	)	,
(	1608	)	,
(	1615	)	,
(	1621	)	,
(	1628	)	,
(	1634	)	,
(	1641	)	,
(	1647	)	,
(	1654	)	,
(	1660	)	,
(	1667	)	,
(	1674	)	,
(	1680	)	,
(	1687	)	,
(	1694	)	,
(	1700	)	,
(	1707	)	,
(	1714	)	,
(	1721	)	,
(	1727	)	,
(	1734	)	,
(	1741	)	,
(	1748	)	,
(	1755	)	,
(	1762	)	,
(	1769	)	,
(	1776	)	,
(	1783	)	,
(	1790	)	,
(	1797	)	,
(	1804	)	,
(	1811	)	,
(	1818	)	,
(	1825	)	,
(	1832	)	,
(	1840	)	,
(	1847	)	,
(	1854	)	,
(	1861	)	,
(	1869	)	,
(	1876	)	,
(	1883	)	,
(	1891	)	,
(	1898	)	,
(	1905	)	,
(	1913	)	,
(	1920	)	,
(	1928	)	,
(	1935	)	,
(	1943	)	,
(	1950	)	,
(	1958	)	,
(	1966	)	,
(	1973	)	,
(	1981	)	,
(	1988	)	,
(	1996	)	,
(	2004	)	,
(	2012	)	,
(	2019	)	,
(	2027	)	,
(	2035	)	,
(	2043	)	,
(	2051	)	,
(	2059	)	,
(	2067	)	,
(	2075	)	,
(	2083	)	,
(	2091	)	,
(	2099	)	,
(	2107	)	,
(	2115	)	,
(	2123	)	,
(	2131	)	,
(	2139	)	,
(	2147	)	,
(	2155	)	,
(	2164	)	,
(	2172	)	,
(	2180	)	,
(	2189	)	,
(	2197	)	,
(	2205	)	,
(	2214	)	,
(	2222	)	,
(	2231	)	,
(	2239	)	,
(	2247	)	,
(	2256	)	,
(	2265	)	,
(	2273	)	,
(	2282	)	,
(	2290	)	,
(	2299	)	,
(	2308	)	,
(	2316	)	,
(	2325	)	,
(	2334	)	,
(	2343	)	,
(	2351	)	,
(	2360	)	,
(	2369	)	,
(	2378	)	,
(	2387	)	,
(	2396	)	,
(	2405	)	,
(	2414	)	,
(	2423	)	,
(	2432	)	,
(	2441	)	,
(	2450	)	,
(	2459	)	,
(	2468	)	,
(	2478	)	,
(	2487	)	,
(	2496	)	,
(	2505	)	,
(	2515	)	,
(	2524	)	,
(	2533	)	,
(	2543	)	,
(	2552	)	,
(	2562	)	,
(	2571	)	,
(	2581	)	,
(	2590	)	,
(	2600	)	,
(	2609	)	,
(	2619	)	,
(	2629	)	,
(	2638	)	,
(	2648	)	,
(	2658	)	,
(	2667	)	,
(	2677	)	,
(	2687	)	,
(	2697	)	,
(	2707	)	,
(	2717	)	,
(	2727	)	,
(	2736	)	,
(	2746	)	,
(	2756	)	,
(	2767	)	,
(	2777	)	,
(	2787	)	,
(	2797	)	,
(	2807	)	,
(	2817	)	,
(	2827	)	,
(	2838	)	,
(	2848	)	,
(	2858	)	,
(	2869	)	,
(	2879	)	,
(	2889	)	,
(	2900	)	,
(	2910	)	,
(	2921	)	,
(	2931	)	,
(	2942	)	,
(	2952	)	,
(	2963	)	,
(	2974	)	,
(	2984	)	,
(	2995	)	,
(	3006	)	,
(	3016	)	,
(	3027	)	,
(	3038	)	,
(	3049	)	,
(	3060	)	,
(	3071	)	,
(	3081	)	,
(	3092	)	,
(	3103	)	,
(	3114	)	,
(	3126	)	,
(	3137	)	,
(	3148	)	,
(	3159	)	,
(	3170	)	,
(	3181	)	,
(	3193	)	,
(	3204	)	,
(	3215	)	,
(	3226	)	,
(	3238	)	,
(	3249	)	,
(	3261	)	,
(	3272	)	,
(	3284	)	,
(	3295	)	,
(	3307	)	,
(	3318	)	,
(	3330	)	,
(	3341	)	,
(	3353	)	,
(	3365	)	,
(	3377	)	,
(	3388	)	,
(	3400	)	,
(	3412	)	,
(	3424	)	,
(	3436	)	,
(	3448	)	,
(	3460	)	,
(	3472	)	,
(	3484	)	,
(	3496	)	,
(	3508	)	,
(	3520	)	,
(	3532	)	,
(	3544	)	,
(	3557	)	,
(	3569	)	,
(	3581	)	,
(	3594	)	,
(	3606	)	,
(	3618	)	,
(	3631	)	,
(	3643	)	,
(	3656	)	,
(	3668	)	,
(	3681	)	,
(	3693	)	,
(	3706	)	,
(	3719	)	,
(	3731	)	,
(	3744	)	,
(	3757	)	,
(	3770	)	,
(	3782	)	,
(	3795	)	,
(	3808	)	,
(	3821	)	,
(	3834	)	,
(	3847	)	,
(	3860	)	,
(	3873	)	,
(	3886	)	,
(	3899	)	,
(	3912	)	,
(	3926	)	,
(	3939	)	,
(	3952	)	,
(	3965	)	,
(	3979	)	,
(	3992	)	,
(	4006	)	,
(	4019	)	,
(	4032	)	,
(	4046	)	,
(	4060	)	,
(	4073	)	,
(	4087	)	,
(	4100	)	,
(	4114	)	,
(	4128	)	,
(	4142	)	,
(	4155	)	,
(	4169	)	,
(	4183	)	,
(	4197	)	,
(	4211	)	,
(	4225	)	,
(	4239	)	,
(	4253	)	,
(	4267	)	,
(	4281	)	,
(	4295	)	,
(	4309	)	,
(	4323	)	,
(	4338	)	,
(	4352	)	,
(	4366	)	,
(	4381	)	,
(	4395	)	,
(	4409	)	,
(	4424	)	,
(	4438	)	,
(	4453	)	,
(	4468	)	,
(	4482	)	,
(	4497	)	,
(	4511	)	,
(	4526	)	,
(	4541	)	,
(	4556	)	,
(	4571	)	,
(	4585	)	,
(	4600	)	,
(	4615	)	,
(	4630	)	,
(	4645	)	,
(	4660	)	,
(	4675	)	,
(	4691	)	,
(	4706	)	,
(	4721	)	,
(	4736	)	,
(	4751	)	,
(	4767	)	,
(	4782	)	,
(	4797	)	,
(	4813	)	,
(	4828	)	,
(	4844	)	,
(	4859	)	,
(	4875	)	,
(	4891	)	,
(	4906	)	,
(	4922	)	,
(	4938	)	,
(	4953	)	,
(	4969	)	,
(	4985	)	,
(	5001	)	,
(	5017	)	,
(	5033	)	,
(	5049	)	,
(	5065	)	,
(	5081	)	,
(	5097	)	,
(	5113	)	,
(	5129	)	,
(	5145	)	,
(	5162	)	,
(	5178	)	,
(	5194	)	,
(	5211	)	,
(	5227	)	,
(	5244	)	,
(	5260	)	,
(	5277	)	,
(	5293	)	,
(	5310	)	,
(	5326	)	,
(	5343	)	,
(	5360	)	,
(	5377	)	,
(	5393	)	,
(	5410	)	,
(	5427	)	,
(	5444	)	,
(	5461	)	,
(	5478	)	,
(	5495	)	,
(	5512	)	,
(	5529	)	,
(	5547	)	,
(	5564	)	,
(	5581	)	,
(	5598	)	,
(	5616	)	,
(	5633	)	,
(	5650	)	,
(	5668	)	,
(	5685	)	,
(	5703	)	,
(	5720	)	,
(	5738	)	,
(	5756	)	,
(	5773	)	,
(	5791	)	,
(	5809	)	,
(	5827	)	,
(	5845	)	,
(	5863	)	,
(	5880	)	,
(	5898	)	,
(	5916	)	,
(	5935	)	,
(	5953	)	,
(	5971	)	,
(	5989	)	,
(	6007	)	,
(	6026	)	,
(	6044	)	,
(	6062	)	,
(	6081	)	,
(	6099	)	,
(	6118	)	,
(	6136	)	,
(	6155	)	,
(	6173	)	,
(	6192	)	,
(	6211	)	,
(	6229	)	,
(	6248	)	,
(	6267	)	,
(	6286	)	,
(	6305	)	,
(	6324	)	,
(	6343	)	,
(	6362	)	,
(	6381	)	,
(	6400	)	,
(	6419	)	,
(	6438	)	,
(	6458	)	,
(	6477	)	,
(	6496	)	,
(	6516	)	,
(	6535	)	,
(	6554	)	,
(	6574	)	,
(	6594	)	,
(	6613	)	,
(	6633	)	,
(	6652	)	,
(	6672	)	,
(	6692	)	,
(	6712	)	,
(	6732	)	,
(	6752	)	,
(	6771	)	,
(	6791	)	,
(	6812	)	,
(	6832	)	,
(	6852	)	,
(	6872	)	,
(	6892	)	,
(	6912	)	,
(	6933	)	,
(	6953	)	,
(	6973	)	,
(	6994	)	,
(	7014	)	,
(	7035	)	,
(	7055	)	,
(	7076	)	,
(	7097	)	,
(	7117	)	,
(	7138	)	,
(	7159	)	,
(	7180	)	,
(	7201	)	,
(	7222	)	,
(	7243	)	,
(	7264	)	,
(	7285	)	,
(	7306	)	,
(	7327	)	,
(	7348	)	,
(	7369	)	,
(	7391	)	,
(	7412	)	,
(	7434	)	,
(	7455	)	,
(	7476	)	,
(	7498	)	,
(	7520	)	,
(	7541	)	,
(	7563	)	,
(	7585	)	,
(	7606	)	,
(	7628	)	,
(	7650	)	,
(	7672	)	,
(	7694	)	,
(	7716	)	,
(	7738	)	,
(	7760	)	,
(	7782	)	,
(	7804	)	,
(	7827	)	,
(	7849	)	,
(	7871	)	,
(	7893	)	,
(	7916	)	,
(	7938	)	,
(	7961	)	,
(	7983	)	,
(	8006	)	,
(	8029	)	,
(	8051	)	,
(	8074	)	,
(	8097	)	,
(	8120	)	,
(	8143	)	,
(	8166	)	,
(	8189	)	,
(	8212	)	,
(	8235	)	,
(	8258	)	,
(	8281	)	,
(	8304	)	,
(	8328	)	,
(	8351	)	,
(	8374	)	,
(	8398	)	,
(	8421	)	,
(	8445	)	,
(	8468	)	,
(	8492	)	,
(	8516	)	,
(	8539	)	,
(	8563	)	,
(	8587	)	,
(	8611	)	,
(	8635	)	,
(	8659	)	,
(	8683	)	,
(	8707	)	,
(	8731	)	,
(	8755	)	,
(	8779	)	,
(	8804	)	,
(	8828	)	,
(	8852	)	,
(	8877	)	,
(	8901	)	,
(	8926	)	,
(	8950	)	,
(	8975	)	,
(	9000	)	,
(	9024	)	,
(	9049	)	,
(	9074	)	,
(	9099	)	,
(	9124	)	,
(	9149	)	,
(	9174	)	,
(	9199	)	,
(	9224	)	,
(	9249	)	,
(	9274	)	,
(	9300	)	,
(	9325	)	,
(	9350	)	,
(	9376	)	,
(	9401	)	,
(	9427	)	,
(	9452	)	,
(	9478	)	,
(	9504	)	,
(	9530	)	,
(	9555	)	,
(	9581	)	,
(	9607	)	,
(	9633	)	,
(	9659	)	,
(	9685	)	,
(	9711	)	,
(	9737	)	,
(	9764	)	,
(	9790	)	,
(	9816	)	,
(	9843	)	,
(	9869	)	,
(	9895	)	,
(	9922	)	,
(	9949	)	,
(	9975	)	,
(	10002	)	,
(	10029	)	,
(	10055	)	,
(	10082	)	,
(	10109	)	,
(	10136	)	,
(	10163	)	,
(	10190	)	,
(	10217	)	,
(	10244	)	,
(	10272	)	,
(	10299	)	,
(	10326	)	,
(	10354	)	,
(	10381	)	,
(	10409	)	,
(	10436	)	,
(	10464	)	,
(	10491	)	,
(	10519	)	,
(	10547	)	,
(	10575	)	,
(	10603	)	,
(	10630	)	,
(	10658	)	,
(	10686	)	,
(	10715	)	,
(	10743	)	,
(	10771	)	,
(	10799	)	,
(	10827	)	,
(	10856	)	,
(	10884	)	,
(	10913	)	,
(	10941	)	,
(	10970	)	,
(	10998	)	,
(	11027	)	,
(	11056	)	,
(	11085	)	,
(	11114	)	,
(	11142	)	,
(	11171	)	,
(	11200	)	,
(	11230	)	,
(	11259	)	,
(	11288	)	,
(	11317	)	,
(	11346	)	,
(	11376	)	,
(	11405	)	,
(	11435	)	,
(	11464	)	,
(	11494	)	,
(	11523	)	,
(	11553	)	,
(	11583	)	,
(	11613	)	,
(	11643	)	,
(	11673	)	,
(	11703	)	,
(	11733	)	,
(	11763	)	,
(	11793	)	,
(	11823	)	,
(	11853	)	,
(	11884	)	,
(	11914	)	,
(	11945	)	,
(	11975	)	,
(	12006	)	,
(	12036	)	,
(	12067	)	,
(	12098	)	,
(	12128	)	,
(	12159	)	,
(	12190	)	,
(	12221	)	,
(	12252	)	,
(	12283	)	,
(	12314	)	,
(	12346	)	,
(	12377	)	,
(	12408	)	,
(	12440	)	,
(	12471	)	,
(	12502	)	,
(	12534	)	,
(	12566	)	,
(	12597	)	,
(	12629	)	,
(	12661	)	,
(	12693	)	,
(	12725	)	,
(	12757	)	,
(	12789	)	,
(	12821	)	,
(	12853	)	,
(	12885	)	,
(	12917	)	,
(	12950	)	,
(	12982	)	,
(	13014	)	,
(	13047	)	,
(	13080	)	,
(	13112	)	,
(	13145	)	,
(	13178	)	,
(	13210	)	,
(	13243	)	,
(	13276	)	,
(	13309	)	,
(	13342	)	,
(	13375	)	,
(	13409	)	,
(	13442	)	,
(	13475	)	,
(	13508	)	,
(	13542	)	,
(	13575	)	,
(	13609	)	,
(	13642	)	,
(	13676	)	,
(	13710	)	,
(	13744	)	,
(	13777	)	,
(	13811	)	,
(	13845	)	,
(	13879	)	,
(	13913	)	,
(	13948	)	,
(	13982	)	,
(	14016	)	,
(	14050	)	,
(	14085	)	,
(	14119	)	,
(	14154	)	,
(	14188	)	,
(	14223	)	,
(	14258	)	,
(	14293	)	,
(	14327	)	,
(	14362	)	,
(	14397	)	,
(	14432	)	,
(	14467	)	,
(	14503	)	,
(	14538	)	,
(	14573	)	,
(	14608	)	,
(	14644	)	,
(	14679	)	,
(	14715	)	,
(	14750	)	,
(	14786	)	,
(	14822	)	,
(	14858	)	,
(	14893	)	,
(	14929	)	,
(	14965	)	,
(	15001	)	,
(	15038	)	,
(	15074	)	,
(	15110	)	,
(	15146	)	,
(	15183	)	,
(	15219	)	,
(	15256	)	,
(	15292	)	,
(	15329	)	,
(	15365	)	,
(	15402	)	,
(	15439	)	,
(	15476	)	,
(	15513	)	,
(	15550	)	,
(	15587	)	,
(	15624	)	,
(	15661	)	,
(	15699	)	,
(	15736	)	,
(	15773	)	,
(	15811	)	,
(	15848	)	,
(	15886	)	,
(	15924	)	,
(	15961	)	,
(	15999	)	,
(	16037	)	,
(	16075	)	,
(	16113	)	,
(	16151	)	,
(	16189	)	,
(	16227	)	,
(	16266	)	,
(	16304	)	,
(	16342	)	,
(	16381	)	,
(	16419	)	,
(	16458	)	,
(	16497	)	,
(	16535	)	,
(	16574	)	,
(	16613	)	,
(	16652	)	,
(	16691	)	,
(	16730	)	,
(	16769	)	,
(	16809	)	,
(	16848	)	,
(	16887	)	,
(	16927	)	,
(	16966	)	,
(	17006	)	,
(	17045	)	,
(	17085	)	,
(	17125	)	,
(	17165	)	,
(	17204	)	,
(	17244	)	,
(	17284	)	,
(	17325	)	,
(	17365	)	,
(	17405	)	,
(	17445	)	,
(	17486	)	,
(	17526	)	,
(	17567	)	,
(	17607	)	,
(	17648	)	,
(	17689	)	,
(	17729	)	,
(	17770	)	,
(	17811	)	,
(	17852	)	,
(	17893	)	,
(	17934	)	,
(	17976	)	,
(	18017	)	,
(	18058	)	,
(	18100	)	,
(	18141	)	,
(	18183	)	,
(	18224	)	,
(	18266	)	,
(	18308	)	,
(	18350	)	,
(	18391	)	,
(	18433	)	,
(	18476	)	,
(	18518	)	,
(	18560	)	,
(	18602	)	,
(	18644	)	,
(	18687	)	,
(	18729	)	,
(	18772	)	,
(	18815	)	,
(	18857	)	,
(	18900	)	,
(	18943	)	,
(	18986	)	,
(	19029	)	,
(	19072	)	,
(	19115	)	,
(	19158	)	,
(	19201	)	,
(	19245	)	,
(	19288	)	,
(	19332	)	,
(	19375	)	,
(	19419	)	,
(	19463	)	,
(	19506	)	,
(	19550	)	,
(	19594	)	,
(	19638	)	,
(	19682	)	,
(	19726	)	,
(	19770	)	,
(	19815	)	,
(	19859	)	,
(	19904	)	,
(	19948	)	,
(	19993	)	,
(	20037	)	,
(	20082	)	,
(	20127	)	,
(	20172	)	,
(	20217	)	,
(	20262	)	,
(	20307	)	,
(	20352	)	,
(	20397	)	,
(	20443	)	,
(	20488	)	,
(	20533	)	,
(	20579	)	,
(	20625	)	,
(	20670	)	,
(	20716	)	,
(	20762	)	,
(	20808	)	,
(	20854	)	,
(	20900	)	,
(	20946	)	,
(	20992	)	,
(	21039	)	,
(	21085	)	,
(	21131	)	,
(	21178	)	,
(	21225	)	,
(	21271	)	,
(	21318	)	,
(	21365	)	,
(	21412	)	,
(	21459	)	,
(	21506	)	,
(	21553	)	,
(	21600	)	,
(	21647	)	,
(	21695	)	,
(	21742	)	,
(	21790	)	,
(	21837	)	,
(	21885	)	,
(	21933	)	,
(	21980	)	,
(	22028	)	,
(	22076	)	,
(	22124	)	,
(	22173	)	,
(	22221	)	,
(	22269	)	,
(	22317	)	,
(	22366	)	,
(	22414	)	,
(	22463	)	,
(	22512	)	,
(	22560	)	,
(	22609	)	,
(	22658	)	,
(	22707	)	,
(	22756	)	,
(	22805	)	,
(	22855	)	,
(	22904	)	,
(	22953	)	,
(	23003	)	,
(	23052	)	,
(	23102	)	,
(	23151	)	,
(	23201	)	,
(	23251	)	,
(	23301	)	,
(	23351	)	,
(	23401	)	,
(	23451	)	,
(	23502	)	,
(	23552	)	,
(	23602	)	,
(	23653	)	,
(	23703	)	,
(	23754	)	,
(	23805	)	,
(	23856	)	,
(	23906	)	,
(	23957	)	,
(	24008	)	,
(	24060	)	,
(	24111	)	,
(	24162	)	,
(	24213	)	,
(	24265	)	,
(	24316	)	,
(	24368	)	,
(	24420	)	,
(	24471	)	,
(	24523	)	,
(	24575	)	,
(	24627	)	,
(	24679	)	,
(	24732	)	,
(	24784	)	,
(	24836	)	,
(	24889	)	,
(	24941	)	,
(	24994	)	,
(	25046	)	,
(	25099	)	,
(	25152	)	,
(	25205	)	,
(	25258	)	,
(	25311	)	,
(	25364	)	,
(	25417	)	,
(	25471	)	,
(	25524	)	,
(	25578	)	,
(	25631	)	,
(	25685	)	,
(	25739	)	,
(	25792	)	,
(	25846	)	,
(	25900	)	,
(	25954	)	,
(	26009	)	,
(	26063	)	,
(	26117	)	,
(	26172	)	,
(	26226	)	,
(	26281	)	,
(	26335	)	,
(	26390	)	,
(	26445	)	,
(	26500	)	,
(	26555	)	,
(	26610	)	,
(	26665	)	,
(	26720	)	,
(	26776	)	,
(	26831	)	,
(	26887	)	,
(	26942	)	,
(	26998	)	,
(	27054	)	,
(	27109	)	,
(	27165	)	,
(	27221	)	,
(	27277	)	,
(	27334	)	,
(	27390	)	,
(	27446	)	,
(	27503	)	,
(	27559	)	,
(	27616	)	,
(	27673	)	,
(	27729	)	,
(	27786	)	,
(	27843	)	,
(	27900	)	,
(	27957	)	,
(	28015	)	,
(	28072	)	,
(	28129	)	,
(	28187	)	,
(	28244	)	,
(	28302	)	,
(	28360	)	,
(	28418	)	,
(	28475	)	,
(	28533	)	,
(	28592	)	,
(	28650	)	,
(	28708	)	,
(	28766	)	,
(	28825	)	,
(	28883	)	,
(	28942	)	,
(	29001	)	,
(	29059	)	,
(	29118	)	,
(	29177	)	,
(	29236	)	,
(	29295	)	,
(	29355	)	,
(	29414	)	,
(	29473	)	,
(	29533	)	,
(	29593	)	,
(	29652	)	,
(	29712	)	,
(	29772	)	,
(	29832	)	,
(	29892	)	,
(	29952	)	,
(	30012	)	,
(	30072	)	,
(	30133	)	,
(	30193	)	,
(	30254	)	,
(	30315	)	,
(	30375	)	,
(	30436	)	,
(	30497	)	,
(	30558	)	,
(	30619	)	,
(	30680	)	,
(	30742	)	,
(	30803	)	,
(	30865	)	,
(	30926	)	,
(	30988	)	,
(	31049	)	,
(	31111	)	,
(	31173	)	,
(	31235	)	,
(	31297	)	,
(	31360	)	,
(	31422	)	,
(	31484	)	,
(	31547	)	,
(	31609	)	,
(	31672	)	,
(	31735	)	,
(	31798	)	,
(	31860	)	,
(	31924	)	,
(	31987	)	,
(	32050	)	,
(	32113	)	,
(	32177	)	,
(	32240	)	,
(	32304	)	,
(	32367	)	,
(	32431	)	,
(	32495	)	,
(	32559	)	,
(	32623	)	,
(	32687	)	,
(	32751	)	,
(	32816	)	,
(	32880	)	,
(	32945	)	,
(	33009	)	,
(	33074	)	,
(	33139	)	,
(	33204	)	,
(	33268	)	,
(	33334	)	,
(	33399	)	,
(	33464	)	,
(	33529	)	,
(	33595	)	,
(	33660	)	,
(	33726	)	,
(	33792	)	,
(	33858	)	,
(	33923	)	,
(	33989	)	,
(	34056	)	,
(	34122	)	,
(	34188	)	,
(	34255	)	,
(	34321	)	,
(	34388	)	,
(	34454	)	,
(	34521	)	,
(	34588	)	,
(	34655	)	,
(	34722	)	,
(	34789	)	,
(	34856	)	,
(	34924	)	,
(	34991	)	,
(	35059	)	,
(	35126	)	,
(	35194	)	,
(	35262	)	,
(	35330	)	,
(	35398	)	,
(	35466	)	,
(	35534	)	,
(	35603	)	,
(	35671	)	,
(	35740	)	,
(	35808	)	,
(	35877	)	,
(	35946	)	,
(	36015	)	,
(	36084	)	,
(	36153	)	,
(	36222	)	,
(	36291	)	,
(	36361	)	,
(	36430	)	,
(	36500	)	,
(	36569	)	,
(	36639	)	,
(	36709	)	,
(	36779	)	,
(	36849	)	,
(	36919	)	,
(	36990	)	,
(	37060	)	,
(	37131	)	,
(	37201	)	,
(	37272	)	,
(	37343	)	,
(	37413	)	,
(	37484	)	,
(	37556	)	,
(	37627	)	,
(	37698	)	,
(	37769	)	,
(	37841	)	,
(	37912	)	,
(	37984	)	,
(	38056	)	,
(	38128	)	,
(	38200	)	,
(	38272	)	,
(	38344	)	,
(	38416	)	,
(	38489	)	,
(	38561	)	,
(	38634	)	,
(	38706	)	,
(	38779	)	,
(	38852	)	,
(	38925	)	,
(	38998	)	,
(	39071	)	,
(	39145	)	,
(	39218	)	,
(	39292	)	,
(	39365	)	,
(	39439	)	,
(	39513	)	,
(	39587	)	,
(	39661	)	,
(	39735	)	,
(	39809	)	,
(	39883	)	,
(	39958	)	,
(	40032	)	,
(	40107	)	,
(	40182	)	,
(	40256	)	,
(	40331	)	,
(	40406	)	,
(	40481	)	,
(	40557	)	,
(	40632	)	,
(	40708	)	,
(	40783	)	,
(	40859	)	,
(	40935	)	,
(	41010	)	,
(	41086	)	,
(	41162	)	,
(	41239	)	,
(	41315	)	,
(	41391	)	,
(	41468	)	,
(	41544	)	,
(	41621	)	,
(	41698	)	,
(	41775	)	,
(	41852	)	,
(	41929	)	,
(	42006	)	,
(	42083	)	,
(	42161	)	,
(	42238	)	,
(	42316	)	,
(	42394	)	,
(	42472	)	,
(	42550	)	,
(	42628	)	,
(	42706	)	,
(	42784	)	,
(	42863	)	,
(	42941	)	,
(	43020	)	,
(	43098	)	,
(	43177	)	,
(	43256	)	,
(	43335	)	,
(	43414	)	,
(	43494	)	,
(	43573	)	,
(	43652	)	,
(	43732	)	,
(	43812	)	,
(	43891	)	,
(	43971	)	,
(	44051	)	,
(	44131	)	,
(	44212	)	,
(	44292	)	,
(	44372	)	,
(	44453	)	,
(	44533	)	,
(	44614	)	,
(	44695	)	,
(	44776	)	,
(	44857	)	,
(	44938	)	,
(	45020	)	,
(	45101	)	,
(	45182	)	,
(	45264	)	,
(	45346	)	,
(	45428	)	,
(	45510	)	,
(	45592	)	,
(	45674	)	,
(	45756	)	,
(	45838	)	,
(	45921	)	,
(	46004	)	,
(	46086	)	,
(	46169	)	,
(	46252	)	,
(	46335	)	,
(	46418	)	,
(	46501	)	,
(	46585	)	,
(	46668	)	,
(	46752	)	,
(	46836	)	,
(	46919	)	,
(	47003	)	,
(	47087	)	,
(	47172	)	,
(	47256	)	,
(	47340	)	,
(	47425	)	,
(	47509	)	,
(	47594	)	,
(	47679	)	,
(	47764	)	,
(	47849	)	,
(	47934	)	,
(	48019	)	,
(	48105	)	,
(	48190	)	,
(	48276	)	,
(	48361	)	,
(	48447	)	,
(	48533	)	,
(	48619	)	,
(	48705	)	,
(	48792	)	,
(	48878	)	,
(	48965	)	,
(	49051	)	,
(	49138	)	,
(	49225	)	,
(	49312	)	,
(	49399	)	,
(	49486	)	,
(	49573	)	,
(	49661	)	,
(	49748	)	,
(	49836	)	,
(	49924	)	,
(	50012	)	,
(	50100	)	,
(	50188	)	,
(	50276	)	,
(	50364	)	,
(	50453	)	,
(	50541	)	,
(	50630	)	,
(	50719	)	,
(	50808	)	,
(	50897	)	,
(	50986	)	,
(	51075	)	,
(	51165	)	,
(	51254	)	,
(	51344	)	,
(	51433	)	,
(	51523	)	,
(	51613	)	,
(	51703	)	,
(	51793	)	,
(	51884	)	,
(	51974	)	,
(	52065	)	,
(	52155	)	,
(	52246	)	,
(	52337	)	,
(	52428	)	,
(	52519	)	,
(	52610	)	,
(	52702	)	,
(	52793	)	,
(	52885	)	,
(	52977	)	,
(	53068	)	,
(	53160	)	,
(	53252	)	,
(	53345	)	,
(	53437	)	,
(	53529	)	,
(	53622	)	,
(	53714	)	,
(	53807	)	,
(	53900	)	,
(	53993	)	,
(	54086	)	,
(	54179	)	,
(	54273	)	,
(	54366	)	,
(	54460	)	,
(	54554	)	,
(	54648	)	,
(	54741	)	,
(	54836	)	,
(	54930	)	,
(	55024	)	,
(	55119	)	,
(	55213	)	,
(	55308	)	,
(	55403	)	,
(	55498	)	,
(	55593	)	,
(	55688	)	,
(	55783	)	,
(	55878	)	,
(	55974	)	,
(	56070	)	,
(	56165	)	,
(	56261	)	,
(	56357	)	,
(	56453	)	,
(	56550	)	,
(	56646	)	,
(	56743	)	,
(	56839	)	,
(	56936	)	,
(	57033	)	,
(	57130	)	,
(	57227	)	,
(	57324	)	,
(	57421	)	,
(	57519	)	,
(	57617	)	,
(	57714	)	,
(	57812	)	,
(	57910	)	,
(	58008	)	,
(	58106	)	,
(	58205	)	,
(	58303	)	,
(	58402	)	,
(	58500	)	,
(	58599	)	,
(	58698	)	,
(	58797	)	,
(	58897	)	,
(	58996	)	,
(	59095	)	,
(	59195	)	,
(	59295	)	,
(	59394	)	,
(	59494	)	,
(	59594	)	,
(	59695	)	,
(	59795	)	,
(	59895	)	,
(	59996	)	,
(	60097	)	,
(	60198	)	,
(	60298	)	,
(	60400	)	,
(	60501	)	,
(	60602	)	,
(	60704	)	,
(	60805	)	,
(	60907	)	,
(	61009	)	,
(	61111	)	,
(	61213	)	,
(	61315	)	,
(	61417	)	,
(	61520	)	,
(	61622	)	,
(	61725	)	,
(	61828	)	,
(	61931	)	,
(	62034	)	,
(	62137	)	,
(	62240	)	,
(	62344	)	,
(	62448	)	,
(	62551	)	,
(	62655	)	,
(	62759	)	,
(	62863	)	,
(	62967	)	,
(	63072	)	,
(	63176	)	,
(	63281	)	,
(	63386	)	,
(	63491	)	,
(	63596	)	,
(	63701	)	,
(	63806	)	,
(	63911	)	,
(	64017	)	,
(	64123	)	,
(	64228	)	,
(	64334	)	,
(	64440	)	,
(	64547	)	,
(	64653	)	,
(	64759	)	,
(	64866	)	,
(	64973	)	,
(	65079	)	,
(	65186	)	,
(	65293	)	,
(	65401	)	,
(	65508	)	,
(	65615	)	,
(	65723	)	,
(	65831	)	,
(	65939	)	,
(	66047	)	,
(	66155	)	,
(	66263	)	,
(	66371	)	,
(	66480	)	,
(	66589	)	,
(	66697	)	,
(	66806	)	,
(	66915	)	,
(	67025	)	,
(	67134	)	,
(	67243	)	,
(	67353	)	,
(	67463	)	,
(	67572	)	,
(	67682	)	,
(	67793	)	,
(	67903	)	,
(	68013	)	,
(	68124	)	,
(	68234	)	,
(	68345	)	,
(	68456	)	,
(	68567	)	,
(	68678	)	,
(	68790	)	,
(	68901	)	,
(	69013	)	,
(	69124	)	,
(	69236	)	,
(	69348	)	,
(	69460	)	,
(	69572	)	,
(	69685	)	,
(	69797	)	,
(	69910	)	,
(	70023	)	,
(	70136	)	,
(	70249	)	,
(	70362	)	,
(	70475	)	,
(	70589	)	,
(	70702	)	,
(	70816	)	,
(	70930	)	,
(	71044	)	,
(	71158	)	,
(	71272	)	,
(	71387	)	,
(	71501	)	,
(	71616	)	,
(	71731	)	,
(	71846	)	,
(	71961	)	,
(	72076	)	,
(	72192	)	,
(	72307	)	,
(	72423	)	,
(	72539	)	,
(	72654	)	,
(	72770	)	,
(	72887	)	,
(	73003	)	,
(	73119	)	,
(	73236	)	,
(	73353	)	,
(	73470	)	,
(	73587	)	,
(	73704	)	,
(	73821	)	,
(	73939	)	,
(	74056	)	,
(	74174	)	,
(	74292	)	,
(	74410	)	,
(	74528	)	,
(	74646	)	,
(	74765	)	,
(	74883	)	,
(	75002	)	,
(	75121	)	,
(	75240	)	,
(	75359	)	,
(	75478	)	,
(	75597	)	,
(	75717	)	,
(	75837	)	,
(	75956	)	,
(	76076	)	,
(	76196	)	,
(	76317	)	,
(	76437	)	,
(	76557	)	,
(	76678	)	,
(	76799	)	,
(	76920	)	,
(	77041	)	,
(	77162	)	,
(	77283	)	,
(	77405	)	,
(	77527	)	,
(	77648	)	,
(	77770	)	,
(	77892	)	,
(	78015	)	,
(	78137	)	,
(	78259	)	,
(	78382	)	,
(	78505	)	,
(	78628	)	,
(	78751	)	,
(	78874	)	,
(	78997	)	,
(	79121	)	,
(	79245	)	,
(	79368	)	,
(	79492	)	,
(	79616	)	,
(	79740	)	,
(	79865	)	,
(	79989	)	,
(	80114	)	,
(	80239	)	,
(	80364	)	,
(	80489	)	,
(	80614	)	,
(	80739	)	,
(	80865	)	,
(	80990	)	,
(	81116	)	,
(	81242	)	,
(	81368	)	,
(	81495	)	,
(	81621	)	,
(	81747	)	,
(	81874	)	,
(	82001	)	,
(	82128	)	,
(	82255	)	,
(	82382	)	,
(	82510	)	,
(	82637	)	,
(	82765	)	,
(	82893	)	,
(	83021	)	,
(	83149	)	,
(	83277	)	,
(	83406	)	,
(	83534	)	,
(	83663	)	,
(	83792	)	,
(	83921	)	,
(	84050	)	,
(	84179	)	,
(	84309	)	,
(	84438	)	,
(	84568	)	,
(	84698	)	,
(	84828	)	,
(	84958	)	,
(	85088	)	,
(	85219	)	,
(	85350	)	,
(	85480	)	,
(	85611	)	,
(	85742	)	,
(	85874	)	,
(	86005	)	,
(	86137	)	,
(	86268	)	,
(	86400	)	,
(	86532	)	,
(	86664	)	,
(	86796	)	,
(	86929	)	,
(	87061	)	,
(	87194	)	,
(	87327	)	,
(	87460	)	,
(	87593	)	,
(	87727	)	,
(	87860	)	,
(	87994	)	,
(	88127	)	,
(	88261	)	,
(	88395	)	,
(	88530	)	,
(	88664	)	,
(	88799	)	,
(	88933	)
);



end package LUT_pkg;
