library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is


type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	4098	)	,
(	4084	)	,
(	4069	)	,
(	4055	)	,
(	4041	)	,
(	4027	)	,
(	4013	)	,
(	3999	)	,
(	3986	)	,
(	3972	)	,
(	3958	)	,
(	3945	)	,
(	3932	)	,
(	3918	)	,
(	3905	)	,
(	3892	)	,
(	3879	)	,
(	3866	)	,
(	3853	)	,
(	3840	)	,
(	3828	)	,
(	3815	)	,
(	3802	)	,
(	3790	)	,
(	3778	)	,
(	3765	)	,
(	3753	)	,
(	3741	)	,
(	3729	)	,
(	3717	)	,
(	3705	)	,
(	3693	)	,
(	3681	)	,
(	3670	)	,
(	3658	)	,
(	3646	)	,
(	3635	)	,
(	3623	)	,
(	3612	)	,
(	3601	)	,
(	3590	)	,
(	3578	)	,
(	3567	)	,
(	3556	)	,
(	3545	)	,
(	3534	)	,
(	3524	)	,
(	3513	)	,
(	3502	)	,
(	3492	)	,
(	3481	)	,
(	3470	)	,
(	3460	)	,
(	3450	)	,
(	3439	)	,
(	3429	)	,
(	3419	)	,
(	3409	)	,
(	3399	)	,
(	3389	)	,
(	3379	)	,
(	3369	)	,
(	3359	)	,
(	3349	)	,
(	3339	)	,
(	3330	)	,
(	3320	)	,
(	3310	)	,
(	3301	)	,
(	3291	)	,
(	3282	)	,
(	3272	)	,
(	3263	)	,
(	3254	)	,
(	3245	)	,
(	3235	)	,
(	3226	)	,
(	3217	)	,
(	3208	)	,
(	3199	)	,
(	3190	)	,
(	3181	)	,
(	3173	)	,
(	3164	)	,
(	3155	)	,
(	3146	)	,
(	3138	)	,
(	3129	)	,
(	3121	)	,
(	3112	)	,
(	3104	)	,
(	3095	)	,
(	3087	)	,
(	3078	)	,
(	3070	)	,
(	3062	)	,
(	3054	)	,
(	3045	)	,
(	3037	)	,
(	3029	)	,
(	3021	)	,
(	3013	)	,
(	3005	)	,
(	2997	)	,
(	2989	)	,
(	2982	)	,
(	2974	)	,
(	2966	)	,
(	2958	)	,
(	2951	)	,
(	2943	)	,
(	2935	)	,
(	2928	)	,
(	2920	)	,
(	2913	)	,
(	2905	)	,
(	2898	)	,
(	2891	)	,
(	2883	)	,
(	2876	)	,
(	2869	)	,
(	2861	)	,
(	2854	)	,
(	2847	)	,
(	2840	)	,
(	2833	)	,
(	2826	)	,
(	2819	)	,
(	2812	)	,
(	2805	)	,
(	2798	)	,
(	2791	)	,
(	2784	)	,
(	2777	)	,
(	2770	)	,
(	2764	)	,
(	2757	)	,
(	2750	)	,
(	2744	)	,
(	2737	)	,
(	2730	)	,
(	2724	)	,
(	2717	)	,
(	2711	)	,
(	2704	)	,
(	2698	)	,
(	2691	)	,
(	2685	)	,
(	2679	)	,
(	2672	)	,
(	2666	)	,
(	2660	)	,
(	2653	)	,
(	2647	)	,
(	2641	)	,
(	2635	)	,
(	2629	)	,
(	2622	)	,
(	2616	)	,
(	2610	)	,
(	2604	)	,
(	2598	)	,
(	2592	)	,
(	2586	)	,
(	2580	)	,
(	2575	)	,
(	2569	)	,
(	2563	)	,
(	2557	)	,
(	2551	)	,
(	2545	)	,
(	2540	)	,
(	2534	)	,
(	2528	)	,
(	2523	)	,
(	2517	)	,
(	2511	)	,
(	2506	)	,
(	2500	)	,
(	2495	)	,
(	2489	)	,
(	2484	)	,
(	2478	)	,
(	2473	)	,
(	2467	)	,
(	2462	)	,
(	2456	)	,
(	2451	)	,
(	2446	)	,
(	2440	)	,
(	2435	)	,
(	2430	)	,
(	2424	)	,
(	2419	)	,
(	2414	)	,
(	2409	)	,
(	2404	)	,
(	2399	)	,
(	2393	)	,
(	2388	)	,
(	2383	)	,
(	2378	)	,
(	2373	)	,
(	2368	)	,
(	2363	)	,
(	2358	)	,
(	2353	)	,
(	2348	)	,
(	2343	)	,
(	2338	)	,
(	2333	)	,
(	2329	)	,
(	2324	)	,
(	2319	)	,
(	2314	)	,
(	2309	)	,
(	2305	)	,
(	2300	)	,
(	2295	)	,
(	2290	)	,
(	2286	)	,
(	2281	)	,
(	2276	)	,
(	2272	)	,
(	2267	)	,
(	2263	)	,
(	2258	)	,
(	2253	)	,
(	2249	)	,
(	2244	)	,
(	2240	)	,
(	2235	)	,
(	2231	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2213	)	,
(	2209	)	,
(	2204	)	,
(	2200	)	,
(	2196	)	,
(	2191	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2174	)	,
(	2170	)	,
(	2166	)	,
(	2162	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2133	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2100	)	,
(	2096	)	,
(	2092	)	,
(	2088	)	,
(	2084	)	,
(	2081	)	,
(	2077	)	,
(	2073	)	,
(	2069	)	,
(	2065	)	,
(	2061	)	,
(	2057	)	,
(	2054	)	,
(	2050	)	,
(	2046	)	,
(	2042	)	,
(	2038	)	,
(	2035	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2020	)	,
(	2016	)	,
(	2013	)	,
(	2009	)	,
(	2005	)	,
(	2002	)	,
(	1998	)	,
(	1994	)	,
(	1991	)	,
(	1987	)	,
(	1984	)	,
(	1980	)	,
(	1977	)	,
(	1973	)	,
(	1970	)	,
(	1966	)	,
(	1963	)	,
(	1959	)	,
(	1956	)	,
(	1952	)	,
(	1949	)	,
(	1945	)	,
(	1942	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1928	)	,
(	1925	)	,
(	1922	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1857	)	,
(	1854	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1820	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1747	)	,
(	1745	)	,
(	1742	)	,
(	1739	)	,
(	1736	)	,
(	1734	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1723	)	,
(	1720	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1709	)	,
(	1707	)	,
(	1704	)	,
(	1701	)	,
(	1699	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1688	)	,
(	1685	)	,
(	1683	)	,
(	1680	)	,
(	1678	)	,
(	1675	)	,
(	1673	)	,
(	1670	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1647	)	,
(	1645	)	,
(	1642	)	,
(	1640	)	,
(	1637	)	,
(	1635	)	,
(	1633	)	,
(	1630	)	,
(	1628	)	,
(	1625	)	,
(	1623	)	,
(	1620	)	,
(	1618	)	,
(	1616	)	,
(	1613	)	,
(	1611	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1597	)	,
(	1594	)	,
(	1592	)	,
(	1590	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1544	)	,
(	1542	)	,
(	1540	)	,
(	1538	)	,
(	1536	)	,
(	1534	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1363	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1318	)	,
(	1317	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	



);



end package LUT_pkg;
